`timescale 1ns / 1ps
module GAME_INTERFACE(clk_25M,hcount,vcount,red,green,blue);
input clk_25M;
input [9:0] hcount,vcount;
output [3:0] red,green,blue;
wire clk_25M;
wire [9:0] hcount,vcount;

wire [0:423] title;
wire [5:0] title_adrs;
wire [0:299] list;
wire [7:0] list_adrs;
wire [0:127] names;
wire [5:0] names_adrs;

Title_Interface Bitmapping_Data(clk_25M,title,title_adrs,list,list_adrs,names,names_adrs);
DISP_WRITE_INTERFACE DISP(clk_25M,hcount,vcount,red,green,blue,title_adrs,title,list,list_adrs,names,names_adrs);

endmodule

module DISP_WRITE_INTERFACE(clk_25M,hcount,vcount,red,green,blue,title_adrs,title,list,list_adrs,names,names_adrs);
input clk_25M;
input [9:0] hcount,vcount;
input [0:423] title;
input [0:299] list;
input [0:127] names;
output reg [5:0] names_adrs;
output reg [7:0] list_adrs;
output reg [5:0] title_adrs;
output reg [3:0] red,green,blue;
always @(posedge clk_25M)
begin
    if((hcount>=144 && hcount<=784) && (vcount>=35 && vcount<=521))
        begin
            title_adrs<=vcount-60;
            list_adrs<=vcount-170;
            names_adrs<=vcount-437;
            if((hcount>252 && hcount<676)&& (vcount>=60 && vcount<115)&& title[hcount-252]==1)
            begin
                {red,green,blue}<={4'b1101,4'b0000,4'b0111};
            end
            else if((hcount>300 && hcount<600)&& (vcount>=170 && vcount<363)&& list[hcount-300]==0)
            begin
                {red,green,blue}<={4'b1101,4'b1100,4'b0111};
            end
            else if((hcount>647 && hcount<775)&& (vcount>=437 && vcount<500)&& names[hcount-647]==1)
            begin
                {red,green,blue}<={4'b1101,4'b1010,4'b1101};
            end
            else
            {red,green,blue}<={4'b0011,4'b0101,4'b0110}; 
        end
    else
        begin
            {red,green,blue}<={4'b0000,4'b0000,4'b0000};   
        end
end
endmodule

module Title_Interface(clk_25M,title,title_adrs,list,list_adrs,names,names_adrs);
input clk_25M;
output reg [0:423] title;
output reg [0:299] list;
output reg [0:127] names;
input [5:0] names_adrs;
input [7:0] list_adrs;
input [5:0] title_adrs;
always @(posedge clk_25M)
begin
    case(title_adrs)
        6'd00:title<=424'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd01:title<=424'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd02:title<=424'b011111111111111111000000000011111111100001111111110000000001111111111000111111111111111111111110000011111111000000000000000000000000000000111111111111111110000000000111111110000000000000000000000000111111111000000011111111100000000000111111111000000001111111111111000000000001111111111111111111100000000000000001111111111110000000000000111111110000000001111111110000011111111100000000011111111000000111111111111111110000000;
6'd03:title<=424'b011111111111111111110000000011111111100000111111111000000001111111110000111111111111111111111110000011111111000000000000000000000000000000111111111111111111100000000111111110000000000000000000000001111111111000000001111111110000000001111111111000000011111111111111100000000001111111111111111111110000000000000011111111111111100000000000111111110000000001111111110000011111111100000000011111111000000111111111111111111000000;
6'd04:title<=424'b011111111111111111111000000011111111100000111111111000000001111111110000111111111111111111111110000011111111000000000000000000000000000000111111111111111111110000000111111110000000000000000000000001111111111100000001111111110000000001111111110000000111111111111111110000000001111111111111111111111000000000000111111111111111110000000000111111110000000001111111110000011111111100000000011111111000000111111111111111111110000;
6'd05:title<=424'b011111111111111111111000000011111111100000111111111000000011111111110000111111111111111111111110000011111111000000000000000000000000000000111111111111111111110000000111111110000000000000000000000001111111111100000001111111110000000001111111110000001111111111111111111000000001111111111111111111111100000000001111111111111111110000000000111111110000000001111111110000011111111110000000011111111000000111111111111111111110000;
6'd06:title<=424'b011111111111111111111100000011111111100000011111111100000011111111100000111111111111111111111110000011111111000000000000000000000000000000111111111111111111111000000111111110000000000000000000000001111111111100000000111111111000000001111111110000011111111111111111111100000001111111111111111111111100000000001111111111111111111000000000111111110000000001111111110000011111111110000000011111111000000111111111111111111111000;
6'd07:title<=424'b011111111111111111111100000011111111100000011111111100000011111111100000111111111111111111111110000011111111000000000000000000000000000000111111111111111111111000000111111110000000000000000000000001111111111100000000111111111000000011111111100000011111111111111111111100000001111111111111111111111110000000011111111111111111111100000000111111110000000001111111110000011111111110000000011111111000000111111111111111111111100;
6'd08:title<=424'b011111111111111111111110000011111111100000011111111100000011111111000000111111111111111111111110000011111111000000000000000000000000000000111111111111111111111100000111111110000000000000000000000011111111111100000000111111111000000011111111100000111111111111111111111100000001111111111111111111111110000000111111111111111111111100000000111111110000000001111111110000011111111111000000011111111000000111111111111111111111100;
6'd09:title<=424'b011111111111111111111110000011111111100000001111111110000111111111000000111111111111111111111110000011111111000000000000000000000000000000111111111111111111111100000111111110000000000000000000000011111111111110000000011111111100000011111111100000111111111111111111111110000001111111111111111111111110000000111111111111111111111110000000111111110000000001111111110000011111111111000000011111111000000111111111111111111111110;
6'd10:title<=424'b011111111111111111111110000011111111100000001111111110000111111111000000111111111111111111111110000011111111000000000000000000000000000000111111111111111111111100000111111110000000000000000000000011111111111110000000011111111100000111111111000001111111111111111111111110000001111111111111111111111111000000111111111111111111111110000000111111110000000001111111110000011111111111100000011111111000000111111111111111111111110;
6'd11:title<=424'b011111111111111111111110000011111111100000001111111110000111111110000000111111111111111111111110000011111111000000000000000000000000000000111111111111111111111100000111111110000000000000000000000011111111111110000000011111111100000111111111000001111111111111111111111110000001111111111111111111111111000001111111111111111111111110000000111111110000000001111111110000011111111111100000011111111000000111111111111111111111110;
6'd12:title<=424'b011111111000001111111110000011111111100000000111111111001111111110000000111111111000000000000000000011111111000000000000000000000000000000111111110000011111111100000111111110000000000000000000000011111111111110000000001111111110000111111110000001111111111000011111111111000001111111110000001111111111000001111111111111111111111111000000111111110000000001111111110000011111111111100000011111111000000111111111111111111111110;
6'd13:title<=424'b011111111000000111111110000011111111100000000111111111001111111110000000111111111000000000000000000011111111000000000000000000000000000000111111110000001111111100000111111110000000000000000000000111111111111110000000001111111110001111111110000011111111110000001111111111000001111111110000000111111111000001111111111000001111111111000000111111110000000001111111110000011111111111110000011111111000000111111111000011111111111;
6'd14:title<=424'b011111111000000111111111000011111111100000000111111111001111111100000000111111111000000000000000000011111111000000000000000000000000000000111111110000001111111100000111111110000000000000000000000111111111111111000000001111111110001111111110000011111111100000000111111111000001111111110000000111111111000011111111110000001111111111000000111111110000000001111111110000011111111111110000011111111000000111111110000001111111111;
6'd15:title<=424'b011111111000000111111111000011111111100000000011111111111111111100000000111111111000000000000000000011111111000000000000000000000000000000111111110000001111111110000111111110000000000000000000000111111111111111000000000111111111001111111100000011111111100000000111111110000001111111110000000111111111000011111111100000000111111111000000111111110000000001111111110000011111111111110000011111111000000111111110000000111111111;
6'd16:title<=424'b011111111000000111111111000011111111100000000011111111111111111100000000111111111000000000000000000011111111000000000000000000000000000000111111110000001111111110000111111110000000000000000000000111111111111111000000000111111111011111111100000011111111000000000011110000000001111111110000000011111111000011111111100000000011111111000000111111110000000001111111110000011111111111111000011111111000000111111110000000111111111;
6'd17:title<=424'b011111111000000111111111000011111111100000000011111111111111111000000000111111111000000000000000000011111111000000000000000000000000000000111111110000001111111110000111111110000000000000000000000111111101111111000000000011111111011111111100000111111111000000000010000000000001111111110000000111111111000011111111100000000011111111100000111111110000000001111111110000011111111111111000011111111000000111111110000000011111111;
6'd18:title<=424'b011111111000000111111111000011111111100000000001111111111111111000000000111111111000000000000000000011111111000000000000000000000000000000111111110000001111111110000111111110000000000000000000001111111101111111000000000011111111111111111000000111111111000000000000000000000001111111110000000111111111000011111111000000000011111111100000111111110000000001111111110000011111111111111000011111111000000111111110000000011111111;
6'd19:title<=424'b011111111000000111111111000011111111100000000001111111111111111000000000111111111000000000000000000011111111000000000000000000000000000000111111110000001111111110000111111110000000000000000000001111111001111111100000000011111111111111111000000111111111000000000000000000000001111111110000000111111111000011111111000000000011111111100000111111110000000001111111110000011111111111111100011111111000000111111110000000011111111;
6'd20:title<=424'b011111111000000111111111000011111111100000000000111111111111110000000000111111111111111111111000000011111111000000000000000000000000000000111111110000001111111100000111111110000000000000000000001111111001111111100000000001111111111111111000000111111111000000000000000000000001111111110000000111111111000111111111000000000001111111100000111111110000000001111111110000011111111111111100011111111000000111111110000000011111111;
6'd21:title<=424'b011111111000000111111110000011111111100000000000111111111111110000000000111111111111111111111100000011111111000000000000000000000000000000111111110000001111111100000111111110000000000000000000001111111001111111100000000001111111111111110000000111111110000000000000000000000001111111110000011111111110000111111111000000000001111111100000111111110000000001111111110000011111111111111110011111111000000111111110000000011111111;
6'd22:title<=424'b011111111000001111111110000011111111100000000000111111111111110000000000111111111111111111111100000011111111000000000000000000000000000000111111110000011111111100000111111110000000000000000000001111111000111111100000000001111111111111110000000111111110000000000000000000000001111111111111111111111110000111111111000000000001111111100000111111110000000001111111110000011111111111111110011111111000000111111110000000011111111;
6'd23:title<=424'b011111111111111111111110000011111111100000000000011111111111100000000000111111111111111111111100000011111111000000000000000000000000000000111111111111111111111100000111111110000000000000000000011111111000111111100000000000111111111111110000000111111110000000111111111111000001111111111111111111111110000111111111000000000001111111100000111111110000000001111111110000011111111111111110011111111000000111111110000000001111111;
6'd24:title<=424'b011111111111111111111110000011111111100000000000011111111111100000000000111111111111111111111100000011111111000000000000000000000000000000111111111111111111111100000111111110000000000000000000011111111000111111110000000000111111111111100000000111111110000001111111111111000001111111111111111111111100000111111111000000000001111111100000111111110000000001111111110000011111111111111111011111111000000111111110000000001111111;
6'd25:title<=424'b011111111111111111111110000011111111100000000000011111111111100000000000111111111111111111111100000011111111000000000000000000000000000000111111111111111111111100000111111110000000000000000000011111111000111111110000000000111111111111100000000111111110000001111111111111000001111111111111111111111100000111111111000000000001111111100000111111110000000001111111110000011111111111111111011111111000000111111110000000001111111;
6'd26:title<=424'b011111111111111111111100000011111111100000000000011111111111100000000000111111111111111111111100000011111111000000000000000000000000000000111111111111111111111000000111111110000000000000000000011111110000111111110000000000011111111111000000000111111110000001111111111111000001111111111111111111111000000111111111000000000001111111100000111111110000000001111111110000011111111111111111011111111000000111111110000000001111111;
6'd27:title<=424'b011111111111111111111100000011111111100000000000011111111111100000000000111111111111111111111100000011111111000000000000000000000000000000111111111111111111111000000111111110000000000000000000011111110000111111110000000000011111111111000000000111111110000001111111111111000001111111111111111111111000000111111111000000000001111111100000111111110000000001111111110000011111111011111111111111111000000111111110000000001111111;
6'd28:title<=424'b011111111111111111111100000011111111100000000000011111111111100000000000111111111111111111111100000011111111000000000000000000000000000000111111111111111111110000000111111110000000000000000000111111110000111111110000000000011111111111000000000111111110000001111111111111000001111111111111111111110000000111111111000000000001111111100000111111110000000001111111110000011111111001111111111111111000000111111110000000001111111;
6'd29:title<=424'b011111111111111111111000000011111111100000000000111111111111110000000000111111111111111111111100000011111111000000000000000000000000000000111111111111111111110000000111111110000000000000000000111111110000011111111000000000001111111110000000000111111110000001111111111111000001111111111111111111000000000111111111000000000001111111100000111111110000000001111111110000011111111001111111111111111000000111111110000000001111111;
6'd30:title<=424'b011111111111111111110000000011111111100000000000111111111111110000000000111111111111111111111100000011111111000000000000000000000000000000111111111111111111100000000111111110000000000000000000111111110000011111111000000000001111111110000000000111111110000001111111111111000001111111111111111111000000000111111111000000000001111111100000111111110000000001111111110000011111111001111111111111111000000111111110000000001111111;
6'd31:title<=424'b011111111111111111100000000011111111100000000001111111111111110000000000111111111000000000000000000011111111000000000000000000000000000000111111111111111111000000000111111110000000000000000000111111110000011111111000000000001111111110000000000111111110000001111111111111000001111111111111111111100000000111111111000000000001111111100000111111110000000001111111110000011111111000111111111111111000000111111110000000001111111;
6'd32:title<=424'b011111111111111111000000000011111111100000000001111111111111111000000000111111111000000000000000000011111111000000000000000000000000000000111111111111111110000000000111111110000000000000000000111111100000011111111000000000001111111110000000000111111110000001111111111111000001111111110011111111110000000111111111000000000001111111100000111111110000000001111111110000011111111000111111111111111000000111111110000000011111111;
6'd33:title<=424'b011111111111100000000000000011111111100000000001111111111111111000000000111111111000000000000000000011111111000000000000000000000000000000111111111111000000000000000111111110000000000000000001111111111111111111111000000000001111111110000000000111111111000000111111111111000001111111110001111111111000000111111111000000000001111111100000111111110000000001111111110000011111111000011111111111111000000111111110000000011111111;
6'd34:title<=424'b011111111000000000000000000011111111100000000011111111111111111000000000111111111000000000000000000011111111000000000000000000000000000000111111110000000000000000000111111110000000000000000001111111111111111111111100000000001111111110000000000111111111000000000001111111000001111111110001111111111000000011111111000000000011111111100000111111110000000001111111110000011111111000011111111111111000000111111110000000011111111;
6'd35:title<=424'b011111111000000000000000000011111111100000000011111111111111111100000000111111111000000000000000000011111111000000000000000000000000000000111111110000000000000000000111111110000000000000000001111111111111111111111100000000001111111110000000000111111111000000000001111111000001111111110000111111111000000011111111000000000011111111100000111111110000000001111111110000011111111000011111111111111000000111111110000000011111111;
6'd36:title<=424'b011111111000000000000000000011111111100000000011111111111111111100000000111111111000000000000000000011111111000000000000000000000000000000111111110000000000000000000111111110000000000000000001111111111111111111111100000000001111111110000000000111111111000000000001111111000001111111110000111111111100000011111111100000000011111111100000111111111000000001111111110000011111111000001111111111111000000111111110000000011111111;
6'd37:title<=424'b011111111000000000000000000011111111100000000111111111011111111100000000111111111000000000000000000011111111000000000000000000000000000000111111110000000000000000000111111110000000000000000001111111111111111111111100000000001111111110000000000011111111000000000001111111000001111111110000111111111100000011111111100000000011111111000000111111111000000001111111100000011111111000001111111111111000000111111110000000111111111;
6'd38:title<=424'b011111111000000000000000000011111111100000000111111111001111111110000000111111111000000000000000000011111111000000000000000000000000000000111111110000000000000000000111111110000000000000000011111111111111111111111100000000001111111110000000000011111111100000000001111111000001111111110000011111111100000011111111100000000111111111000000111111111000000011111111100000011111111000001111111111111000000111111110000000111111111;
6'd39:title<=424'b011111111000000000000000000011111111100000000111111111001111111110000000111111111000000000000000000011111111000000000000000000000000000000111111110000000000000000000111111111000000000000000011111111111111111111111110000000001111111110000000000011111111100000000011111111000001111111110000011111111110000011111111110000000111111111000000111111111100000011111111100000011111111000000111111111111000000111111110000001111111111;
6'd40:title<=424'b011111111000000000000000000011111111100000001111111110001111111110000000111111111000000000000000000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111100011111111111111111111111110000000001111111110000000000011111111110000000111111111000001111111110000011111111110000001111111111000001111111111000000011111111110000111111111100000011111111000000111111111111000000111111111000011111111111;
6'd41:title<=424'b011111111000000000000000000011111111100000001111111110000111111111000000111111111111111111111110000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111100011111111111111111111111110000000001111111110000000000001111111111000001111111111000001111111110000001111111110000001111111111111111111111111000000011111111111111111111111100000011111111000000111111111111000000111111111111111111111111;
6'd42:title<=424'b011111111000000000000000000011111111100000001111111110000111111111000000111111111111111111111110000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111100011111111111111111111111110000000001111111110000000000001111111111111111111111111000001111111110000001111111110000001111111111111111111111110000000011111111111111111111111100000011111111000000011111111111000000111111111111111111111110;
6'd43:title<=424'b011111111000000000000000000011111111100000011111111100000111111111100000111111111111111111111110000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111100111111111111111111111111110000000001111111110000000000001111111111111111111111111000001111111110000001111111111000000111111111111111111111110000000011111111111111111111111000000011111111000000011111111111000000111111111111111111111110;
6'd44:title<=424'b011111111000000000000000000011111111100000011111111100000011111111100000111111111111111111111110000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111100111111110000000000111111111000000001111111110000000000000111111111111111111111111000001111111110000001111111111000000111111111111111111111100000000001111111111111111111111000000011111111000000001111111111000000111111111111111111111100;
6'd45:title<=424'b011111111000000000000000000011111111100000111111111100000011111111100000111111111111111111111110000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111100111111110000000000111111111000000001111111110000000000000111111111111111111111111000001111111110000000111111111000000111111111111111111111100000000001111111111111111111111000000011111111000000001111111111000000111111111111111111111100;
6'd46:title<=424'b011111111000000000000000000011111111100000111111111000000011111111110000111111111111111111111110000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111100111111110000000000111111111000000001111111110000000000000011111111111111111111110000001111111110000000111111111100000011111111111111111111100000000001111111111111111111110000000011111111000000001111111111000000111111111111111111111000;
6'd47:title<=424'b011111111000000000000000000011111111100000111111111000000001111111110000111111111111111111111110000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111100111111110000000000011111111000000001111111110000000000000011111111111111111111100000001111111110000000111111111100000001111111111111111111000000000000111111111111111111110000000011111111000000000111111111000000111111111111111111111000;
6'd48:title<=424'b011111111000000000000000000011111111100001111111111000000001111111110000111111111111111111111110000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111101111111110000000000011111111000000001111111110000000000000001111111111111111111000000001111111110000000011111111100000001111111111111111110000000000000011111111111111111100000000011111111000000000111111111000000111111111111111111110000;
6'd49:title<=424'b011111111000000000000000000011111111100001111111110000000001111111111000111111111111111111111110000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111101111111110000000000011111111100000001111111110000000000000000111111111111111110000000001111111110000000011111111100000000111111111111111100000000000000011111111111111111000000000011111111000000000111111111000000111111111111111111100000;
6'd50:title<=424'b011111111000000000000000000011111111100001111111110000000000111111111000111111111111111111111110000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111101111111100000000000011111111100000001111111110000000000000000011111111111111100000000001111111110000000011111111110000000011111111111111100000000000000001111111111111110000000000011111111000000000011111111000000111111111111111111000000;
6'd51:title<=424'b011111111000000000000000000011111111100011111111110000000000111111111000111111111111111111111110000011111111111111111111100000000000000000111111110000000000000000000111111111111111111111101111111100000000000011111111100000001111111110000000000000000001111111111111000000000001111111110000000011111111110000000001111111111110000000000000000000111111111111100000000000011111111000000000011111111000000111111111111111100000000;
6'd52:title<=424'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000;
6'd53:title<=424'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd54:title<=424'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        default: title<=0;
    endcase
end

always @(list_adrs)
begin
    case(list_adrs)
    8'd000:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd001:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd002:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd003:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd004:list<=300'b111111111111111111100001111111111111111000000000000011111111000011110000011111111000011111111000000000011111111111111111111100000000001111111111111000001111111111000000011111110000001111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd005:list<=300'b111111111111111111100001111111111111111000000000000001111111000011110000011111111000011111110000000000001111111111111111111000000000000111111111111000001111111111000000011111110000001111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd006:list<=300'b111111111111111111000001111111111111111000000000000000111111000011110000001111111000011111100000000000000111111111111111110000000000000011111111111000000111111111000000011111100000001111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd007:list<=300'b111111111111111111000001111111111111111000000000000000111111000011110000001111111000011111000000000000000011111111111111100000000000000011111111111000000111111111000000011111100000001111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd008:list<=300'b111111111111111110000001111111111111111000001110000000011111000011110000001111111000011111000000111100000011111111111111100000011110000001111111110000000111111111000000011111100000001111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd009:list<=300'b111111111111111100000001111111111111111000001111110000011111000011110000000111111000011110000001111110000001111111111111000001111111000001111111110000000011111111000000001111100000001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd010:list<=300'b111111111111111000000001111111111111111000001111111000001111000011110000000111111000011110000011111111000001111111111111000011111111100001111111110000000011111111000000001111100000001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd011:list<=300'b111111111111110000000001111111111111111000001111111100001111000011110000000011111000011110000111111111100001111111111110000011111111100001111111100000000011111111000000001111100000001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd012:list<=300'b111111111111110000000001111111111111111000001111111100001111000011110000000011111000011110000111111111100001111111111110000011111111100111111111100001000011111111000000001111000000001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd013:list<=300'b111111111111110000100001111111111111111000001111111100001111000011110000000001111000011100000111111111100000111111111110000111111111111111111111100001000001111111000010001111000000001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd014:list<=300'b111111111111110001100001111111111111111000001111111100000111000011110000000001111000011100000111111111100000111111111110000111111111111111111111100001100001111111000010000111000100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd015:list<=300'b111111111111110011100001111111111111111000001111111100000111000011110000100001111000011100001111111111110000111111111110000111111111111111111111000011100001111111000010000111000100001111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd016:list<=300'b111111111111111111100001111111111111111000001111111100000111000011110000100000111000011100001111111111110000111111111110000111111111111111111111000011100000111111000010000111000100001111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd017:list<=300'b111111111111111111100001111111111111111000001111111100000111000011110000110000111000011100001111111111110000111111111110000111111000000001111111000011110000111111000011000110000100001111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd018:list<=300'b111111111111111111100001111111111111111000001111111100000111000011110000110000011000011100001111111111110000111111111110000111111000000000111110000011110000111111000011000110000100001111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd019:list<=300'b111111111111111111100001111111111111111000001111111100000111000011110000111000011000011100001111111111110000111111111110000111111000000000111110000111110000111111000011000010000100001111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd020:list<=300'b111111111111111111100001111111111111111000001111111100000111000011110000111000001000011100001111111111110000111111111110000111111000000000111110000111110000011111000011000010001100001111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd021:list<=300'b111111111111111111100001111111111111111000001111111100000111000011110000111000001000011100000111111111110000111111111110000111111000000000111110000000000000011111000011000010001100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd022:list<=300'b111111111111111111100001111111111111111000001111111100001111000011110000111100000000011100000111111111100000111111111110000111111111100000111100000000000000011111000011000000001100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd023:list<=300'b111111111111111111100001111111111111111000001111111100001111000011110000111100000000011100000111111111100000111111111110000111111111110000111100000000000000001111000011100000001100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd024:list<=300'b111111111111111111100001111111111111111000001111111100001111000011110000111110000000011110000111111111100001111111111110000011111111110000111100000000000000001111000011100000001100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd025:list<=300'b111111111111111111100001111111111111111000001111111000001111000011110000111110000000011110000011111111000001111111111111000011111111110000111100000000000000001111000011100000001100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd026:list<=300'b111111111111111111100001111111111111111000001111111000001111000011110000111111000000011110000011111111000001111111111111000001111111100000111000001111111100001111000011100000011100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd027:list<=300'b111111111111111111100001111110000111111000001111110000011111000011110000111111000000011111000001111110000011111111111111000000111111000000111000011111111100000111000011100000011100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd028:list<=300'b111111111111111111100001111110000111111000000000000000011111000011110000111111000000011111000000000000000011111111111111100000000000000000111000011111111100000111000011110000011100001111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd029:list<=300'b111111111111111111100001111110000111111000000000000000111111000011110000111111100000011111100000000000000111111111111111110000000000000001110000011111111110000111000011110000011100001111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd030:list<=300'b111111111111111111100001111110000111111000000000000001111111000011110000111111100000011111110000000000001111111111111111110000000000000011110000011111111110000011000011110000011100001111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd031:list<=300'b111111111111111111100001111110000111111000000000000011111111000011110000111111110000011111111000000000011111111111111111111000000000000111110000111111111110000011000011110000011100001111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd032:list<=300'b111111111111111111100001111110000111111100000000001111111111000011110000111111110000111111111100000000111111111111111111111110000000011111110000111111111111000011000011110000111100001111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd033:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd034:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd035:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd036:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd037:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd038:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd039:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd040:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd041:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd042:list<=300'b111111111111111111000111111111111111110000000000000000111000011111111110000001111111111111111000000000000000011111100001111111111111111100000011111111111111110000000000000000111111100000001111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd043:list<=300'b111111111111111100000001111111111111110000000000000000011000011111111000000000011111111111111000000000000000011111100000111111111111110000000001111111111111100000000000000000111111000000000011111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd044:list<=300'b111111111111111000000000111111111111110000000000000000011000011111110000000000001111111111111000000000000000011111000000111111111111100000000000111111111111100000000000000000111110000000000001111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd045:list<=300'b111111111111110000000000011111111111110000000000000000011000011111100000000000001111111111111000000000000000011111000000111111111111000000000000011111111111100000000000000000111100000000000000111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd046:list<=300'b111111111111100000000000011111111111110000000000000000011000011111000000000000000111111111111000000000000000011111000000011111111110000000000000001111111111100000000000000000111000000000000000111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd047:list<=300'b111111111111100000110000001111111111111111110000011111111000011111000001111100000111111111111111111000011111111111000000011111111110000011111000001111111111111111100000111111111000001111100000011111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd048:list<=300'b111111111111100001111000001111111111111111110000011111111000011111000011111110000011111111111111111000011111111110000000011111111100000111111100000111111111111111110000111111110000011111110000011111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd049:list<=300'b111111111111100001111100001111111111111111110000011111111000011110000011111110000011111111111111111000011111111110000000011111111100000111111100000111111111111111110000111111110000111111111000001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd050:list<=300'b111111111111100001111100001111111111111111110000011111111000011110000111111111000011111111111111111000011111111110000000001111111100001111111110000111111111111111110000111111100000111111111100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd051:list<=300'b111111111111111111111100001111111111111111110000011111111000011110000111111111111111111111111111111000011111111110000100001111111100001111111111111111111111111111110000111111100000111111111100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd052:list<=300'b111111111111111111111100001111111111111111110000011111111000011110000111111111111111111111111111111000011111111100001100001111111000001111111111111111111111111111110000111111100001111111111100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd053:list<=300'b111111111111111111111100001111111111111111110000011111111000011100000111111111111111111111111111111000011111111100001100000111111000001111111111111111111111111111110000111111100001111111111100000111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd054:list<=300'b111111111111111111111000011111111111111111110000011111111000011100000111111111111111111111111111111000011111111100001110000111111000011111111111111111111111111111110000111111100001111111111100000111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd055:list<=300'b111111111111111111111000011111111111111111110000011111111000011100000111111111111111111111111111111000011111111000001110000111111000011111111111111111111111111111110000111111100001111111111100000111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd056:list<=300'b111111111111111111110000111111111111111111110000011111111000011100001111111111111111111111111111111000011111111000011110000111111000011111111111111111111111111111110000111111100001111111111100000111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd057:list<=300'b111111111111111111100000111111111111111111110000011111111000011100000111111111111111111111111111111000011111111000011110000011111000011111111111111111111111111111110000111111100001111111111100000111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd058:list<=300'b111111111111111111000001111111111111111111110000011111111000011100000111111111111111111111111111111000011111111000011111000011111000011111111111111111111111111111110000111111100001111111111100000111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd059:list<=300'b111111111111111111000001111111111111111111110000011111111000011100000111111111111111111111111111111000011111110000011111000011111000001111111111111111111111111111110000111111100001111111111100000111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd060:list<=300'b111111111111111110000011111111111111111111110000011111111000011100000111111111111111111111111111111000011111110000000000000001111000001111111111111111111111111111110000111111100001111111111100000111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd061:list<=300'b111111111111111100000111111111111111111111110000011111111000011110000111111111001111111111111111111000011111110000000000000001111000001111111110011111111111111111110000111111100001111111111100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd062:list<=300'b111111111111111000001111111111111111111111110000011111111000011110000111111111000011111111111111111000011111110000000000000001111100001111111110000111111111111111110000111111100000111111111100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd063:list<=300'b111111111111111000011111111111111111111111110000011111111000011110000111111110000011111111111111111000011111100000000000000001111100001111111100000111111111111111110000111111100000111111111000001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd064:list<=300'b111111111111110000011111111111111111111111110000011111111000011110000011111110000011111111111111111000011111100000000000000000111100000111111100000111111111111111110000111111110000011111111000001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd065:list<=300'b111111111111110000111111111111111111111111110000011111111000011111000001111100000111111111111111111000011111100001111111100000111110000011111000001111111111111111110000111111110000011111110000011111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd066:list<=300'b111111111111100000000000001110000111111111110000011111111000011111000000111000000111111111111111111000011111000001111111110000111110000001110000001111111111111111110000111111111000001111100000011111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd067:list<=300'b111111111111100000000000001110000111111111110000011111111000011111100000000000001111111111111111111000011111000011111111110000011111000000000000011111111111111111110000111111111000000000000000111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd068:list<=300'b111111111111100000000000001110000111111111110000011111111000011111100000000000001111111111111111111000011111000011111111110000011111000000000000011111111111111111110000111111111100000000000000111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd069:list<=300'b111111111111000000000000001110000111111111110000011111111000011111110000000000011111111111111111111000011111000011111111111000011111100000000000111111111111111111110000111111111110000000000001111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd070:list<=300'b111111111111000000000000001110000111111111110000011111111000011111111100000000111111111111111111111000011110000011111111111000011111111000000001111111111111111111110000111111111111000000000011111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd071:list<=300'b111111111111100000000000001110000111111111111000111111111000011111111111000111111111111111111111111000111110000111111111111000011111111110001111111111111111111111110001111111111111110000001111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd072:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd073:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd074:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd075:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd076:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd077:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd078:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd079:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd080:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd081:list<=300'b111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111000000111111111111111100000111111111111111111111111111111111111111111111111;
8'd082:list<=300'b111111111111111100000011111111111111111000000000000011111111111110000000001111111110000000000000111111111111100000111111111100000000000000011110000000111111100000011111111000000000011111111000001111111100001111111111111111100000000001111111111110000000001111111111111111111111111111111111111111111111;
8'd083:list<=300'b111111111111111000000001111111111111111000000000000001111111111000000000000111111110000000000000011111111111100000111111111100000000000000011110000000111111000000011111110000000000001111111100001111111100001111111111111111000000000000111111111100000000000011111111111111111111111111111111111111111111;
8'd084:list<=300'b111111111111110000000000111111111111111000000000000000111111110000000000000011111110000000000000001111111111000000111111111100000000000000011110000000111111000000011111100000000000000111111100000111111100001111111111111110000000000000111111111000000000000001111111111111111111111111111111111111111111;
8'd085:list<=300'b111111111111110000000000011111111111111000000000000000111111110000000000000001111110000000000000000111111111000000011111111100000000000000011110000000111111000000011111100000000000000011111100000111111100001111111111111100000000000000011111110000000000000001111111111111111111111111111111111111111111;
8'd086:list<=300'b111111111111100000000000011111111111111000001111000000011111100000011110000001111110000111111000000111111111000000011111111100000111111111111110000000111111000000011111000000111100000011111100000011111100001111111111111000000111110000001111110000001111000000111111111111111111111111111111111111111111;
8'd087:list<=300'b111111111111100001111000011111111111111000001111110000011111100000111111100000111110000111111100000111111111000000011111111100001111111111111110000000111111000000011111000001111111000001111100000011111100001111111111111000001111111000001111100000111111100000111111111111111111111111111111111111111111;
8'd088:list<=300'b111111111111100001111000011111111111111000001111111000001111000001111111100000111110000111111110000111111110000000001111111100001111111111111110000000011111000000011110000011111111000001111100000001111100001111111111111000011111111100001111100000111111110000011111111111111111111111111111111111111111;
8'd089:list<=300'b111111111111110011111000011111111111111000001111111100001111000001111111110000011110000111111110000111111110000000001111111100001111111111111110000000011110000000011110000011111111100000111100000001111100001111111111110000011111111100001111100001111111110000011111111111111111111111111111111111111111;
8'd090:list<=300'b111111111111111111111000011111111111111000001111111100001111000011111111110000011110000111111110000111111110000100001111111100001111111111111110000000011110000000011110000111111111100000111100000001111100001111111111110000111111111100111111000001111111111000011111111111111111111111111111111111111111;
8'd091:list<=300'b111111111111111111111000011111111111111000001111111100001111000011111111111000011110000111111110000111111110000100001111111100001111111111111110000100011110000000011110000111111111110000111100000000111100001111111111110000111111111111111111000011111111111000011111111111111111111111111111111111111111;
8'd092:list<=300'b111111111111111111110000011111111111111000001111111100000111000011111111111000011110000111111100000111111100001100000111111100001111111111111110000100011110001000011110000111111111110000111100000000111100001111111111110000111111111111111111000011111111111000001111111111111111111111111111111111111111;
8'd093:list<=300'b111111111111111111000000111111111111111000001111111100000110000011111111111000011110000111110000000111111100001110000111111100000000000000111110000100001110001000011100000111111111110000111100010000011100001111111111110000111111111111111111000011111111111000001111111111111111111111111111111111111111;
8'd094:list<=300'b111111111111111111000001111111111111111000001111111100000110000011111111111000011110000000000000001111111100001110000111111100000000000000011110000100001100001000011100000111111111110000111100011000011100001111111111100000111111111111111111000011111111111000001111111111111111111111111111111111111111;
8'd095:list<=300'b111111111111111111000001111111111111111000001111111100000110000011111111111000011110000000000000001111111000001110000011111100000000000000011110000100001100001000011100000111111111110000111100011000001100001111111111100000111111000000001111000011111111111000001111111111111111111111111111111111111111;
8'd096:list<=300'b111111111111111111000000111111111111111000001111111100000110000011111111111000011110000000000000011111111000011110000011111100000000000000011110000110001100001000011100000111111111110000111100011000001100001111111111100000111111000000000111000011111111111000001111111111111111111111111111111111111111;
8'd097:list<=300'b111111111111111111000000011111111111111000001111111100000110000011111111111000011110000000000001111111111000011111000011111100000000000000111110000110001100011000011100000111111111110000111100011100001100001111111111100000111111000000000111000011111111111000001111111111111111111111111111111111111111;
8'd098:list<=300'b111111111111111111111000001111111111111000001111111100000110000011111111111000011110000110000001111111111000011111000011111100001111111111111110000110001100011000011100000111111111110000111100011100000100001111111111110000111111000000000111000011111111111000001111111111111111111111111111111111111111;
8'd099:list<=300'b111111111111111111111100001111111111111000001111111100000110000011111111111000011110000111000000111111110000000000000001111100001111111111111110000110000000011000011100000111111111110000111100011110000100001111111111110000111111000000000111000011111111111000001111111111111111111111111111111111111111;
8'd100:list<=300'b111111111111111111111100001111111111111000001111111100001111000011111111111000011110000111100000111111110000000000000001111100001111111111111110000110000000011000011110000111111111110000111100011110000000001111111111110000111111111100000111000011111111111000011111111111111111111111111111111111111111;
8'd101:list<=300'b111111111111100011111100001111111111111000001111111100001111000001111111110000011110000111110000011111100000000000000000111100001111111111111110000111000000111000011110000011111111100000111100011111000000001111111111110000011111111110000111000001111111111000011111111111111111111111111111111111111111;
8'd102:list<=300'b111111111111100001111100001111111111111000001111111000001111000001111111110000111110000111111000001111100000000000000000111100001111111111111110000111000000111000011110000011111111100001111100011111000000001111111111111000011111111110000111100001111111110000011111111111111111111111111111111111111111;
8'd103:list<=300'b111111111111100001111100001111111111111000001111111000001111100000111111100000111110000111111000001111100001111111100000111100001111111111111110000111000000111000011111000001111111000001111100011111100000001111111111111000001111111100000111100000111111100000111111111111111111111111111111111111111111;
8'd104:list<=300'b111111111111100001111000001110000111111000001111110000011111100000011111000000111110000111111100000111100001111111110000111100001111111111111110000111000000111000011111000000111110000001111100011111100000001111111111111000000111111000000111100000011111000000111111111111111111111111111111111111111111;
8'd105:list<=300'b111111111111100000000000011110000111111000000000000000011111110000000000000001111110000111111100000111000001111111110000011100000000000000001110000111000000111000011111000000000000000011111100011111110000001111111111111100000000000000000111110000000000000000111111111111111111111111111111111111111111;
8'd106:list<=300'b111111111111110000000000011110000111111000000000000000111111110000000000000011111110000111111100000011000011111111110000011100000000000000001110000111000000111000011111100000000000000111111100011111110000001111111111111100000000000000001111111000000000000001111111111111111111111111111111111111111111;
8'd107:list<=300'b111111111111110000000000111110000111111000000000000001111111111000000000000011111110000111111110000011000011111111111000011100000000000000001110000111100001111000011111110000000000000111111100011111111000001111111111111110000000000000011111111000000000000011111111111111111111111111111111111111111111;
8'd108:list<=300'b111111111111111000000001111110000111111000000000000011111111111100000000000111111110000111111110000011000011111111111000001100000000000000001110000111100001111000011111111000000000001111111000011111111000001111111111111111000000000000111111111100000000000111111111111111111111111111111111111111111111;
8'd109:list<=300'b111111111111111100000011111110000111111100000000001111111111111111000000011111111110000111111111000000000011111111111000001100000000000000001110000111100001111000011111111110000000111111111100011111111100001111111111111111110000000011111111111111000000001111111111111111111111111111111111111111111111;
8'd110:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd111:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd112:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd113:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd114:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd115:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd116:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd117:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd118:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd119:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd120:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd121:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd122:list<=300'b111111111111111111111111111111111111111100000000001111111110001111100001111111100001111111111000000011111111111111111100000000001111111111111100000001111111111000011111111100011111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd123:list<=300'b111111111111111111110000111111111111111000000000000011111100000111100001111111100001111111110000000000111111111111111100000000000001111111111000000000011111111000001111111100001111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd124:list<=300'b111111111111111111110000111111111111111000000000000001111100000111100000111111100001111111100000000000011111111111111100000000000000111111110000000000001111111000001111111100001111111000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd125:list<=300'b111111111111111111100000111111111111111000000000000000111100000111100000111111100001111111000000000000001111111111111100000000000000111111100000000000000111111000000111111100001111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd126:list<=300'b111111111111111111100000111111111111111000000000000000111100000111100000111111100001111110000000000000001111111111111100000000000000011111000000000000000011111000000111111100001111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd127:list<=300'b111111111111111111000000111111111111111000001111100000011100000111100000011111100001111100000011111000000111111111111100001111100000011111000001111110000011111000000011111100001111100000011111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd128:list<=300'b111111111111111111000000111111111111111000001111110000011100000111100000011111100001111100000111111100000111111111111100001111110000011110000011111111000001111000000011111100001111100000111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd129:list<=300'b111111111111111111000000111111111111111000001111111000011100000111100000001111100001111100001111111110000111111111111100001111111000011110000011111111000001111000000011111100001111000001111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd130:list<=300'b111111111111111110000000111111111111111000001111111000011100000111100000001111100001111000001111111110000111111111111100001111111000011110000111111111100001111000000001111100001111000011111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd131:list<=300'b111111111111111110000000111111111111111000001111111000011100000111100000000111100001111000011111111111111111111111111100001111111000011100000111111111100001111000000001111100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd132:list<=300'b111111111111111100000000111111111111111000001111111000011100000111100000000111100001111000011111111111111111111111111100001111111000011100000111111111100000111000000000111100001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd133:list<=300'b111111111111111100010000111111111111111000001111111000011100000111100000000111100001111000011111111111111111111111111100001111111000011100001111111111100000111000000000111100001110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd134:list<=300'b111111111111111000010000111111111111111000001111110000011100000111100010000011100001111000011111111111111111111111111100001111110000011100001111111111110000111000010000011100001110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd135:list<=300'b111111111111111000110000111111111111111000001111000000011100000111100011000011100001111000011111111111111111111111111100001111000000011100001111111111110000111000010000011100001110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd136:list<=300'b111111111111110000110000111111111111111000000000000000111100000111100011000001100001111000011111100000000011111111111100000000000000111100001111111111110000111000011000011100001110000011111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd137:list<=300'b111111111111110001110000111111111111111000000000000000111100000111100011100001100001111000011111100000000011111111111100000000000000111100001111111111110000111000011000001100001110000011111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd138:list<=300'b111111111111100001110000111111111111111000000000000001111100000111100011100000100001111000011111100000000011111111111100000000000001111100001111111111110000111000011100001100001110000011111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd139:list<=300'b111111111111100011110000111111111111111000000000000011111100000111100011100000100001111000011111100000000011111111111100000000000011111100001111111111110000111000011100000100001110000011111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd140:list<=300'b111111111111000011110000111111111111111000001111111111111100000111100011110000000001111000011111100000000011111111111100000111111111111100000111111111100000111000011110000000001110000011111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd141:list<=300'b111111111111000000000000000111111111111000001111111111111100000111100011110000000001111000011111111111000011111111111100001111111111111100000111111111100000111000011110000000001111000011111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd142:list<=300'b111111111111000000000000000111111111111000001111111111111100000111100011111000000001111000001111111111000011111111111100001111111111111100000111111111100001111000011110000000001111000011111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd143:list<=300'b111111111111000000000000000111111111111000001111111111111100000111100011111000000001111000001111111111000011111111111100001111111111111110000111111111100001111000011111000000001111000001111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd144:list<=300'b111111111111000000000000000111111111111000001111111111111100000111100011111100000001111100001111111111000011111111111100001111111111111110000011111111000001111000011111000000001111000001111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd145:list<=300'b111111111111000000000000000111111111111000001111111111111100000111100011111100000001111100000111111110000011111111111100001111111111111110000001111110000001111000011111100000001111100000111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd146:list<=300'b111111111111111111110000111110000111111000001111111111111100000111100011111110000001111110000011111000000011111111111100001111111111111111000000111100000011111000011111100000001111100000011111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd147:list<=300'b111111111111111111110000111110000111111000001111111111111100000111100011111110000001111110000000000000000011111111111100001111111111111111000000000000000011111000011111110000001111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd148:list<=300'b111111111111111111110000111110000111111000001111111111111100000111100011111110000001111111000000000000000111111111111100001111111111111111100000000000000111111000011111110000001111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd149:list<=300'b111111111111111111110000111110000111111000001111111111111100000111100011111111000001111111100000000000001111111111111100001111111111111111110000000000001111111000011111110000001111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd150:list<=300'b111111111111111111110000111110000111111000001111111111111100000111100011111111000001111111110000000000111111111111111100001111111111111111111000000000011111111000011111111000001111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd151:list<=300'b111111111111111111111000111110000111111100011111111111111110001111100011111111100011111111111100000011111111111111111100011111111111111111111110000001111111111100011111111100011111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd152:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd153:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd154:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd155:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd156:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd157:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd158:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd159:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd160:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd161:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd162:list<=300'b111111111111111100000000011111111111111000000000000111111111111110000000011111111110000000000011111111111111100000000111111111000000000000000111111111111111110000000111111111111110000011111111110000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd163:list<=300'b111111111111111000000000001111111111111000000000000001111111111100000000000111111110000000000000111111111110000000000011111111000000000000000111111111111111000000000001111111111110000011111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd164:list<=300'b111111111111111000000000001111111111111000000000000000111111111000000000000011111110000000000000011111111100000000000001111111000000000000000111111111111110000000000000111111111110000011111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd165:list<=300'b111111111111111000000000001111111111111000000000000000111111110000000000000001111110000000000000011111111000000000000000111111000000000000000111111111111110000000000000111111111110000001111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd166:list<=300'b111111111111111000000000001111111111111000000000000000011111100000001100000001111110000000000000001111111000000011000000111111000000000000000111111111111100000001000000011111111100000001111111110000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd167:list<=300'b111111111111111000000000001111111111111000001111110000011111100000111111000000111110000111111000001111110000001111110000011111000011111111111111111111111100000111110000011111111100000001111111110000111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd168:list<=300'b111111111111110000111111111111111111111000001111111000001111100000111111100000111110000111111100000111110000011111110000011111000011111111111111111111111000001111111000001111111100000000111111110000111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd169:list<=300'b111111111111110000111111111111111111111000001111111000001111000001111111110000111110000111111100000111110000111111111000011111000011111111111111111111111000011111111000001111111000000000111111110000111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd170:list<=300'b111111111111110000111111111111111111111000001111111100001111000011111111110000011110000111111110000111100000111111111000011111000011111111111111111111111000011111111100011111111000010000111111110000111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd171:list<=300'b111111111111110000111111111111111111111000001111111100001111000011111111111000011110000111111110000111100001111111111111111111000011111111111111111111110000011111111111111111111000010000111111110000111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd172:list<=300'b111111111111110000100011111111111111111000001111111100001111000011111111111000011110000111111110000011100001111111111111111111000011111111111111111111110000011111111111111111111000011000011111110000111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd173:list<=300'b111111111111110000000001111111111111111000001111111100000110000011111111111000011110000111111110000011100001111111111111111111000011111111111111111111110000111111111111111111110000111000011111110000011111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd174:list<=300'b111111111111110000000000111111111111111000001111111100000110000011111111111000011110000111111110000011100001111111111111111111000000000000001111111111110000111111111111111111110000111000011111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd175:list<=300'b111111111111110000000000011111111111111000001111111100000110000011111111111000011110000111111110000011100001111111111111111111000000000000001111111111110000111111111111111111110000111000001111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd176:list<=300'b111111111111100000000000001111111111111000001111111100000110000011111111111000011110000111111110000011100001111110000000001111000000000000001111111111110000111111111111111111100000111100001111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd177:list<=300'b111111111111100000111000001111111111111000001111111100000110000011111111111000011110000111111110000011100001111110000000001111000000000000001111111111110000111111111111111111100001111100001111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd178:list<=300'b111111111111100001111100001111111111111000001111111100000110000011111111111000011110000111111110000011100001111110000000001111000011111111111111111111110000111111111111111111100001111100001111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd179:list<=300'b111111111111111111111100001111111111111000001111111100000110000011111111111000011110000111111110000011100001111110000000001111000011111111111111111111110000111111111111111111100001111100000111110000111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd180:list<=300'b111111111111111111111100001111111111111000001111111100000111000011111111111000011110000111111110000011100001111110000000001111000011111111111111111111110000011111111111111111000000000000000111110000111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd181:list<=300'b111111111111111111111100001111111111111000001111111100001111000011111111111000011110000111111110000111100001111111111100001111000011111111111111111111110000011111111100011111000000000000000111110000111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd182:list<=300'b111111111111111111111100001111111111111000001111111100001111000011111111110000011110000111111110000111100000111111111100001111000011111111111111111111111000011111111000001111000000000000000011110000111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd183:list<=300'b111111111111100001111100001111111111111000001111111100001111000001111111110000011110000111111110000111110000111111111100001111000011111111111111111111111000011111111000001111000000000000000011110000111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd184:list<=300'b111111111111100001111100001111111111111000001111111000001111000001111111100000111110000111111100000111110000011111111000001111000011111111111111111111111000001111111000011110000000000000000011110000111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd185:list<=300'b111111111111100000111100001111111111111000001111110000011111100000111111000000111110000111111000001111110000001111110000001111000011111111111111111111111100000111110000011110000111111111000011110000111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd186:list<=300'b111111111111100000111000001110000111111000000000000000011111100000001110000001111110000000000000001111111000000111100000001111000000000000000111111111111100000000000000011110000111111111000001110000111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd187:list<=300'b111111111111110000000000011110000111111000000000000000111111110000000000000001111110000000000000001111111000000000000000001111000000000000000111111111111110000000000000111100000111111111100001110000111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd188:list<=300'b111111111111110000000000011110000111111000000000000000111111111000000000000011111110000000000000011111111100000000000000011111000000000000000111111111111111000000000001111100000111111111100001110000111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd189:list<=300'b111111111111111000000000111110000111111000000000000001111111111000000000000111111110000000000000111111111110000000000000111111000000000000000111111111111111100000000011111100001111111111100000110000111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd190:list<=300'b111111111111111100000001111110000111111000000000000111111111111110000000001111111110000000000011111111111111000000000011111111000000000000000111111111111111110000000111111100001111111111100000110000111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd191:list<=300'b111111111111111111000111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'd192:list<=300'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    endcase
end
always @(names_adrs)
begin
   case(names_adrs)
   6'd00:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd01:names<=128'b00000000000000000000000000000000000000000000111110000100000110000000000000000000000000000000000000000000000000000000000000000000;
6'd02:names<=128'b00000000000000000000000000000000000000000001111111100110000110000000000000000000000000000000000000000000000000000000000000000000;
6'd03:names<=128'b00000000000000000000000000000000000000000001100001100011001100000000000000000000000000000000000000000000000000000000000000000000;
6'd04:names<=128'b00000000000000000000000000000000000000000001100001100011011000000000000000000000000000000000000000000000000000000000000000000000;
6'd05:names<=128'b00000000000000000000000000000000000000000001111111000001111000000000000000000000000000000000000000000000000000000000000000000000;
6'd06:names<=128'b00000000000000000000000000000000000000000001111111100000110000000000000000000000000000000000000000000000000000000000000000000000;
6'd07:names<=128'b00000000000000000000000000000000000000000001100001100000110000000000000000000000000000000000000000000000000000000000000000000000;
6'd08:names<=128'b00000000000000000000000000000000000000000001100001110000110000000000000000000000000000000000000000000000000000000000000000000000;
6'd09:names<=128'b00000000000000000000000000000000000000000001110011100000110000000000000000000000000000000000000000000000000000000000000000000000;
6'd10:names<=128'b00000000000000000000000000000000000000000001111111100000110000000000000000000000000000000000000000000000000000000000000000000000;
6'd11:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd12:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd13:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd14:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd15:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd16:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd17:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd18:names<=128'b00001110000110000001111111100010000011011000001100000010001100000011001100000110000110011111000001100001000111110000000010000000;
6'd19:names<=128'b00001110001111000001111111100111000011011000001100000111000110001110001100000111000110011111110001100001100111111100000111000000;
6'd20:names<=128'b00001111001111000000001100000011000110011000001100000111000111001100011110000111000110011000111001100001100110001110000111000000;
6'd21:names<=128'b00001111001111000000001100000011000110011000001100001111100011011000011110000111100110011000011001100001100110000110001111100000;
6'd22:names<=128'b00001111011111000000001100000011100110011000001100001101100001111000111011000111100110011000011001111111100111111100001101100000;
6'd23:names<=128'b00001101011011000000001100000001101100011000001100011000110001110000110001000110110110011000011001111111100111111000011000110000;
6'd24:names<=128'b00001101111011000000001100000001101100011000001100011111110000110000111111000110011110011000011001100001100110011000011111110000;
6'd25:names<=128'b00001101110011000000001100000001111100011011001100011111110000110001111111100110011110011000011001100001100110011100011111110000;
6'd26:names<=128'b00001101110011001100001100110000111000011011101100110000011000110001100001100110001110011000110001100001100110001100110000011000;
6'd27:names<=128'b00001100110011001100001100110000111000011001111100110000011000110011000000110110001110011111110001100001100110000110110000011100;
6'd28:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd29:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd30:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd31:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd32:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd33:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd34:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd35:names<=128'b00001111110000000001111000000111100001000011000010011000011100100000110001100000000001110000011111000011000000000000000000000000;
6'd36:names<=128'b00001111111000000011111100001111111001100011100110011100011100110001100011100000000111111100111111110011000000000000000000000000;
6'd37:names<=128'b00001100001100000011000110011100011001100111100110011100111100111001100011110000000110001100110000110011000000000000000000000000;
6'd38:names<=128'b00001100001100000011000000011000001101100111100110011100111100011011000111110000000110000000110000110011000000000000000000000000;
6'd39:names<=128'b00001111111000000011111000011000001100110110100110011110111100001111000110110000000111110000111111110011000000000000000000000000;
6'd40:names<=128'b00001111111000000001111110011000001100110100111100010110101100001110000110011000000001111100111111100011000000000000000000000000;
6'd41:names<=128'b00001100001100000000000110011000001100111100111100010111101100000110001111111000000000001100110011100011000000000000000000000000;
6'd42:names<=128'b00001100001100000110000110011000011100111100111100010011101100000110001111111100000110000110110001100011000000000000000000000000;
6'd43:names<=128'b00001110011100110011001110011100111000011100011100010011101100000110001100001100000111001100110000110011000000000000000000000000;
6'd44:names<=128'b00001111111000110001111100001111110000011000011000010011001100000110011000001100000011111100110000111011000000000000000000000000;
6'd45:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd46:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd47:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd48:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd49:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd50:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd51:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd52:names<=128'b00000001110000110000110000000111100001111110000000100001000000101100000100001000000000000000000000000000000000000000000000000000;
6'd53:names<=128'b00000111111000110000110000001111110001111111000001110001100001101110001100011100000000000000000000000000000000000000000000000000;
6'd54:names<=128'b00001110001100110000110000001100111001100011100001110001100001100110011100011100000000000000000000000000000000000000000000000000;
6'd55:names<=128'b00001100000000110000110000001100000001100001100011111000110001100011011000111110000000000000000000000000000000000000000000000000;
6'd56:names<=128'b00001100000000111111110000001111100001111111000011011000110011000011110000110110000000000000000000000000000000000000000000000000;
6'd57:names<=128'b00001100000000111111110000000111110001111110000011001100111011000001110000110011000000000000000000000000000000000000000000000000;
6'd58:names<=128'b00001100000000110000110000000000111001100110000111111100011011000001100001111111000000000000000000000000000000000000000000000000;
6'd59:names<=128'b00001100001100110000110000001100011001100111000111111110011110000001100001111111000000000000000000000000000000000000000000000000;
6'd60:names<=128'b00000111011100110000110011001100111001100011101110000110011110000001100011000001100000000000000000000000000000000000000000000000;
6'd61:names<=128'b00000011111000110000110011001111110001100001101100000110001110000001100011000001100000000000000000000000000000000000000000000000;
6'd62:names<=128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
   endcase
end
endmodule

