module DORAEMON_GO(sys_clk,clk_25M,clk_100,red,green,blue,hcount,vcount,jump,reset1,rst_dg);
input sys_clk,clk_25M,clk_100,jump,reset1,rst_dg;
output [3:0] red,green,blue;
input [9:0] hcount,vcount;
wire stop,reset,set1;
wire [9:0] hbird=250;
wire [9:0] vbird,obs,entry,obs2,obs3,entry2,entry3;
wire [5:0] data_adrs,go_adrs;
wire [0:39] data;
wire [4:0] score_adrs;
wire [0:19] score1,score2,score3,score4;
wire [3:0] bcd3,bcd2,bcd1,bcd0;
wire [15:0] bcd;
wire [0:99] score_t;
wire [0:235] game_over;
assign bcd3=bcd[15:12];
assign bcd2=bcd[11:8];
assign bcd1=bcd[7:4];
assign bcd0=bcd[3:0];
assign stop_temp=0;
wire reset;
assign reset=reset1|rst_dg;
SCORE_DG Score_counter(sys_clk,bcd,stop,reset);
SCORE_DATA_DG Score1(clk_25M,bcd0,score1,score_adrs,score_t);
SCORE_DATA_DG Score2(clk_25M,bcd1,score2,score_adrs);
SCORE_DATA_DG Score3(clk_25M,bcd2,score3,score_adrs);
SCORE_DATA_DG Score4(clk_25M,bcd3,score4,score_adrs);
DISP_WRITE_DG Disp(clk_25M,hcount,vcount,stop,hbird,vbird,obs,obs2,obs3,entry,entry2,entry3,data_adrs,data,score1,score2,score3,score4,score_t,score_adrs,go_adrs,game_over,red,green,blue);
MOV_BIRD Moving(clk_100,jump,stop,reset,vbird);
OBSTACLE Obstacle(clk_100,jump,obs,obs2,obs3,vbird,hbird,entry,entry2,entry3,stop,reset,set1);
LFSR_FLAPPY LFSR(clk_100,reset,obs,obs2,obs3,entry,entry2,entry3);
DATA_DG DORAEMON(clk_25M,data_adrs,data,go_adrs,game_over);
endmodule

module DISP_WRITE_DG(clk,hcount,vcount,stop,hbird,vbird,obs,obs2,obs3,entry,entry2,entry3,data_adrs,data,score1,score2,score3,score4,score_t,score_adrs,go_adrs,game_over,red,green,blue);
input clk,stop;
input [9:0] hcount,vcount,hbird,vbird,obs,entry,obs2,obs3,entry2,entry3;
output reg [3:0] red,green,blue;
input [0:39] data;
output reg [5:0] data_adrs,go_adrs;
input [0:19] score1;
input [0:19] score2;
input [0:19] score3;
input [0:19] score4;
input [0:99] score_t;
input [0:235] game_over;
output reg [4:0] score_adrs;
always @(posedge clk)
begin
    if((hcount>=144 && hcount<=784) && (vcount>=35 && vcount<=521))
    begin
        data_adrs<=vcount-vbird;
        score_adrs<=vcount-40;
        go_adrs<=vcount-263;
        if((hcount>hbird && hcount<hbird+40)&& (vcount>vbird && vcount<vbird+50) && (data[hcount-hbird]==1))
        begin
            {red,green,blue}={4'b0011,4'b1010,4'b1101};
        end
        else if((hcount>=346 && hcount<=582) && (vcount>=263 && vcount<=327)&&(game_over[hcount-346]==1)&& stop)
            begin
                {red,green,blue}<={4'b1111,4'b0000,4'b0000};
            end
        else if((hcount>=750 && hcount<=770) && (vcount>=40 && vcount<=72)&&(score1[hcount-750]==1))
        begin
            {red,green,blue}<={4'b0000,4'b0000,4'b0000};
        end
        else if((hcount>=730 && hcount<=750) && (vcount>=40 && vcount<=72)&&(score2[hcount-730]==1))
        begin
            {red,green,blue}<={4'b0000,4'b0000,4'b0000};
        end
        else if((hcount>=710 && hcount<=730) && (vcount>=40 && vcount<=72)&&(score3[hcount-710]==1))
        begin
            {red,green,blue}<={4'b0000,4'b0000,4'b0000};
        end
        else if((hcount>=690 && hcount<=710) && (vcount>=40 && vcount<=72)&&(score4[hcount-690]==1))
        begin
            {red,green,blue}<={4'b0000,4'b0000,4'b0000};
        end
        else if((hcount>=590 && hcount<=689) && (vcount>=40 && vcount<=72)&&(score_t[hcount-590]==1))
        begin
            {red,green,blue}<={4'b0000,4'b0000,4'b0000};
        end
        else if(hcount>obs && hcount<=obs+30 && vcount>35 && vcount<=525)
        begin
            if(vcount>entry && vcount <entry+120)
                {red,green,blue}={4'b1111,4'b1111,4'b1101};
            else
                {red,green,blue}={4'b0001,4'b0110,4'b0000};
        end
        else if(hcount>obs2 && hcount<=obs2+30 && vcount>35 && vcount<=525)
        begin
            if(vcount>entry2 && vcount <entry2+120)
                {red,green,blue}={4'b1111,4'b1111,4'b1101};
            else
                {red,green,blue}={4'b0001,4'b0110,4'b0000};
        end
        else if(hcount>obs3 && hcount<=obs3+30 && vcount>35 && vcount<=525)
        begin
            if(vcount>entry3 && vcount <entry3+120)
                {red,green,blue}={4'b1111,4'b1111,4'b1101};
            else
                {red,green,blue}={4'b0001,4'b0110,4'b0000};
        end
        else
        begin
            {red,green,blue}={4'b1111,4'b1111,4'b1101};
        end
    end
    else
    begin
        {red,green,blue}={4'b0000,4'b0000,4'b0000};
    end
end
endmodule

//Obstacle Logic
module OBSTACLE(clk,jump,obs,obs2,obs3,vbird,hbird,entry,entry2,entry3,stop,reset,set1);
input clk,reset,jump;
input [9:0] hbird,vbird,entry,entry2,entry3;
output reg [9:0] obs=500,obs2=800,obs3=100;
output reg stop,set1;
always @(posedge clk)
begin
    if(vbird>=475 || vbird<=35 || ((vbird>entry+70 ||(vbird<=entry-7))&&(obs>hbird-30 && obs<=hbird+35))|| ((vbird>entry2+70 ||(vbird<=entry2-7))&&(obs2>hbird-30 && obs2<=hbird+35))||((vbird>entry3+70 ||(vbird<=entry3-7))&&(obs3>hbird-30 && obs3<=hbird+35)))
    begin
        stop<=1;
    end
    else
        stop<=0;
end
always@(posedge clk)
begin
    if(reset)
    begin
        obs<=500;
        obs2<=800;
        obs3<=77;
        set1<=1;
    end
    else
    begin
        if(stop)
            if(jump)
            begin
                set1<=1;
                obs<=obs;
                obs2<=obs2;
                obs3<=obs3;
            end
            else
            begin
                set1<=0;
                obs<=obs;
                obs2<=obs2;
                obs3<=obs3;
            end
        else
        begin
            obs<=obs-1;
            obs2<=obs2-1;
            obs3<=obs3-1;
            set1<=0;
        end
    end
end
endmodule
// Bird Moving Logic
module MOV_BIRD(clk_10Hz,jump,stop,reset,vbird);
input clk_10Hz,jump,stop,reset;
output reg [9:0] vbird=250;
always @(posedge clk_10Hz)
begin
    if(reset)
        vbird<=250;
    else if(stop)
        vbird<=vbird;
    else if(jump)
        vbird<=vbird-1;
    else
        vbird<=vbird+1;
end
endmodule

// LFSR For Random Obstacles
module LFSR_FLAPPY(clk,reset,obs,obs2,obs3,entry,entry2,entry3);
    input clk,reset;
    input [9:0] obs,obs2,obs3;
    output reg[9:0] entry=50,entry2=200,entry3=300;

    reg [8:0] lfsr;
    wire feedback;

    // Feedback polynomial: x^9 + x^5 + 1
    assign feedback = lfsr[8] ^ lfsr[4];

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            lfsr <= 9'b110010101; // Initialize LFSR to a non-zero value
        end else begin
            lfsr <= {lfsr[7:0], feedback}; // Shift and feedback
        end
    end

    always @(posedge clk) begin
        // Map LFSR output to the range 75 to 360 for different entries
        if(obs<114 || obs> 784)
            entry <= (lfsr % (360 - 75 + 1)) + 75;
        else
            entry<=entry;
        if(obs2<114 || obs2> 784)
            entry2 <= ((lfsr + 123) % (360 - 75 + 1)) + 75; // Offset to generate a different value
        else
            entry2<=entry2;
        if(obs3<114 || obs3> 784)
            entry3 <= ((lfsr + entry-50) % (360 - 75 + 1)) + 75; // Another offset for a unique value
        else
            entry3<=entry3;
    end
endmodule

module SCORE_DG(clk,score,stop_temp,reset);
input clk,reset,stop_temp;
output [15:0] score;
reg clk_div;
integer i;
integer div;
reg [13:0] bin=0;
always @(posedge clk)
begin
    if(i==div)
    begin
        clk_div<=~clk_div;
        i<=0;
    end
    else
        i<=i+1;
end
always @(posedge clk)
begin
    if(bin <15)
        div<=49999999;
    else if( bin>=15 && bin <=30)
        div<=25999999;
    else if( bin>30 && bin <=50)
        div<=12599999;
    else if( bin>50 && bin <=100)
        div<=10000000;
    else if( bin>100 && bin <=1000)
        div<=4999999;
    else if( bin>1000 && bin <10000)
        div<=2599999;
    else
        div<=div;
end
always @(posedge clk_div, posedge reset)
begin
    if(reset)
        bin<=0;
    else if(stop_temp)
        bin<=bin;
    else
        bin<=bin+1;
end
BIN_BCD Binary_BCD(clk,bin,score);
endmodule

module SCORE_DATA_DG(clk_25MHz,count,data,data_adrs,score_t);
input clk_25MHz;
input [4:0] data_adrs;
input [3:0] count;
output reg [0:19] data;
output reg [0:99] score_t;
always @(posedge clk_25MHz)
begin
    case(count)
    4'd0:
        begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000011000000000;
        5'd03:data<=20'b00000011111111000000;
        5'd04:data<=20'b00000111111111100000;
        5'd05:data<=20'b00001111111111110000;
        5'd06:data<=20'b00001111111111110000;
        5'd07:data<=20'b00011111000011111000;
        5'd08:data<=20'b00011110000011111000;
        5'd09:data<=20'b00011110000001111000;
        5'd10:data<=20'b00111110000001111000;
        5'd11:data<=20'b00111110000001111000;
        5'd12:data<=20'b00111110000001111100;
        5'd13:data<=20'b00111100000001111100;
        5'd14:data<=20'b00111100000001111100;
        5'd15:data<=20'b00111100000001111100;
        5'd16:data<=20'b00111100000001111100;
        5'd17:data<=20'b00111100000001111100;
        5'd18:data<=20'b00111100000001111100;
        5'd19:data<=20'b00111110000001111100;
        5'd20:data<=20'b00111110000001111000;
        5'd21:data<=20'b00111110000001111000;
        5'd22:data<=20'b00111110000001111000;
        5'd23:data<=20'b00111110000011111000;
        5'd24:data<=20'b00011111000011111000;
        5'd25:data<=20'b00011111100111110000;
        5'd26:data<=20'b00011111111111110000;
        5'd27:data<=20'b00001111111111100000;
        5'd28:data<=20'b00000111111111000000;
        5'd29:data<=20'b00000011111110000000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;    
        endcase
        end
    4'd1:begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000000000000000;
        5'd04:data<=20'b00000001111000000000;
        5'd05:data<=20'b00000011111000000000;
        5'd06:data<=20'b00000111111000000000;
        5'd07:data<=20'b00011111111000000000;
        5'd08:data<=20'b00011111111000000000;
        5'd09:data<=20'b00011101111000000000;
        5'd10:data<=20'b00011001111000000000;
        5'd11:data<=20'b00000001111000000000;
        5'd12:data<=20'b00000001111000000000;
        5'd13:data<=20'b00000001111000000000;
        5'd14:data<=20'b00000001111000000000;
        5'd15:data<=20'b00000001111000000000;
        5'd16:data<=20'b00000001111000000000;
        5'd17:data<=20'b00000001111000000000;
        5'd18:data<=20'b00000001111000000000;
        5'd19:data<=20'b00000001111000000000;
        5'd20:data<=20'b00000001111000000000;
        5'd21:data<=20'b00000001111000000000;
        5'd22:data<=20'b00000001111000000000;
        5'd23:data<=20'b00000001111000000000;
        5'd24:data<=20'b00000001111000000000;
        5'd25:data<=20'b00000001111100000000;
        5'd26:data<=20'b00011111111111100000;
        5'd27:data<=20'b00011111111111100000;
        5'd28:data<=20'b00011111111111100000;
        5'd29:data<=20'b00011111111111100000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
        end
    4'd2:
        begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000001111100000000;
        5'd03:data<=20'b00000111111111000000;
        5'd04:data<=20'b00011111111111100000;
        5'd05:data<=20'b00011111111111100000;
        5'd06:data<=20'b00011111111111110000;
        5'd07:data<=20'b00011100011111110000;
        5'd08:data<=20'b00011000001111110000;
        5'd09:data<=20'b00000000000111110000;
        5'd10:data<=20'b00000000000111110000;
        5'd11:data<=20'b00000000000111110000;
        5'd12:data<=20'b00000000000111110000;
        5'd13:data<=20'b00000000001111110000;
        5'd14:data<=20'b00000000001111100000;
        5'd15:data<=20'b00000000001111100000;
        5'd16:data<=20'b00000000011111000000;
        5'd17:data<=20'b00000000111111000000;
        5'd18:data<=20'b00000000111110000000;
        5'd19:data<=20'b00000001111100000000;
        5'd20:data<=20'b00000011111000000000;
        5'd21:data<=20'b00000111111000000000;
        5'd22:data<=20'b00001111110000000000;
        5'd23:data<=20'b00001111100000000000;
        5'd24:data<=20'b00011111000000000000;
        5'd25:data<=20'b00011111111111111000;
        5'd26:data<=20'b00111111111111111000;
        5'd27:data<=20'b00111111111111111000;
        5'd28:data<=20'b00011111111111111000;
        5'd29:data<=20'b00011111111111110000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
        end
    4'd3:
        begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000011000000000;
            5'd03:data<=20'b00000111111111000000;
            5'd04:data<=20'b00001111111111100000;
            5'd05:data<=20'b00011111111111100000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011100001111110000;
            5'd08:data<=20'b00010000000111110000;
            5'd09:data<=20'b00000000000111110000;
            5'd10:data<=20'b00000000000111110000;
            5'd11:data<=20'b00000000000111110000;
            5'd12:data<=20'b00000000000111110000;
            5'd13:data<=20'b00000000001111100000;
            5'd14:data<=20'b00000111111111000000;
            5'd15:data<=20'b00001111111110000000;
            5'd16:data<=20'b00001111111111000000;
            5'd17:data<=20'b00000111111111110000;
            5'd18:data<=20'b00000000011111110000;
            5'd19:data<=20'b00000000000111111000;
            5'd20:data<=20'b00000000000011111000;
            5'd21:data<=20'b00000000000011111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011111000;
            5'd24:data<=20'b00010000000111111000;
            5'd25:data<=20'b00111100001111111000;
            5'd26:data<=20'b00111111111111110000;
            5'd27:data<=20'b00111111111111100000;
            5'd28:data<=20'b00011111111111000000;
            5'd29:data<=20'b00001111111110000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
            endcase
        end
    4'd4:
    begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000011111100000;
        5'd04:data<=20'b00000000011111100000;
        5'd05:data<=20'b00000000111111100000;
        5'd06:data<=20'b00000000111111100000;
        5'd07:data<=20'b00000001111111100000;
        5'd08:data<=20'b00000001111111100000;
        5'd09:data<=20'b00000011110111100000;
        5'd10:data<=20'b00000011110111100000;
        5'd11:data<=20'b00000111100111100000;
        5'd12:data<=20'b00000111100111100000;
        5'd13:data<=20'b00001111000111100000;
        5'd14:data<=20'b00001111000111100000;
        5'd15:data<=20'b00011110000111100000;
        5'd16:data<=20'b00011110000111100000;
        5'd17:data<=20'b00111100000111100000;
        5'd18:data<=20'b00111100000111100000;
        5'd19:data<=20'b00111000000111100000;
        5'd20:data<=20'b00111111111111111100;
        5'd21:data<=20'b00111111111111111100;
        5'd22:data<=20'b00111111111111111100;
        5'd23:data<=20'b00111111111111111100;
        5'd24:data<=20'b00000000000111110000;
        5'd25:data<=20'b00000000000111100000;
        5'd26:data<=20'b00000000000111100000;
        5'd27:data<=20'b00000000000111100000;
        5'd28:data<=20'b00000000000111100000;
        5'd29:data<=20'b00000000000111100000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd5:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00001111111111100000;
            5'd04:data<=20'b00011111111111110000;
            5'd05:data<=20'b00011111111111110000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011111111111100000;
            5'd08:data<=20'b00011110000000000000;
            5'd09:data<=20'b00011110000000000000;
            5'd10:data<=20'b00011110000000000000;
            5'd11:data<=20'b00011110000000000000;
            5'd12:data<=20'b00011110000000000000;
            5'd13:data<=20'b00011111111100000000;
            5'd14:data<=20'b00011111111111000000;
            5'd15:data<=20'b00011111111111100000;
            5'd16:data<=20'b00011111111111110000;
            5'd17:data<=20'b00001100011111111000;
            5'd18:data<=20'b00000000000111111000;
            5'd19:data<=20'b00000000000011111000;
            5'd20:data<=20'b00000000000011111000;
            5'd21:data<=20'b00000000000011111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011111000;
            5'd24:data<=20'b00000000000111111000;
            5'd25:data<=20'b00011000001111110000;
            5'd26:data<=20'b00011111111111110000;
            5'd27:data<=20'b00011111111111100000;
            5'd28:data<=20'b00011111111111000000;
            5'd29:data<=20'b00001111111100000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd6:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00000000111111110000;
            5'd04:data<=20'b00000011111111110000;
            5'd05:data<=20'b00000011111111110000;
            5'd06:data<=20'b00000111111111110000;
            5'd07:data<=20'b00001111100000000000;
            5'd08:data<=20'b00001111000000000000;
            5'd09:data<=20'b00011111000000000000;
            5'd10:data<=20'b00011110000000000000;
            5'd11:data<=20'b00011110000000000000;
            5'd12:data<=20'b00011110000000000000;
            5'd13:data<=20'b00011110011111000000;
            5'd14:data<=20'b00011111111111110000;
            5'd15:data<=20'b00011111111111111000;
            5'd16:data<=20'b00111111111111111000;
            5'd17:data<=20'b00111111000011111100;
            5'd18:data<=20'b00111110000001111100;
            5'd19:data<=20'b00011110000001111100;
            5'd20:data<=20'b00011110000001111100;
            5'd21:data<=20'b00011110000001111100;
            5'd22:data<=20'b00011110000001111100;
            5'd23:data<=20'b00011110000001111100;
            5'd24:data<=20'b00011111000001111000;
            5'd25:data<=20'b00011111100011111000;
            5'd26:data<=20'b00001111111111111000;
            5'd27:data<=20'b00001111111111110000;
            5'd28:data<=20'b00000111111111100000;
            5'd29:data<=20'b00000001111110000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd7:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00011111111111111000;
            5'd04:data<=20'b00111111111111111000;
            5'd05:data<=20'b00111111111111111000;
            5'd06:data<=20'b00111111111111111000;
            5'd07:data<=20'b00011111111111111000;
            5'd08:data<=20'b00000000000011111000;
            5'd09:data<=20'b00000000000011111000;
            5'd10:data<=20'b00000000000111110000;
            5'd11:data<=20'b00000000000111110000;
            5'd12:data<=20'b00000000000111110000;
            5'd13:data<=20'b00000000001111100000;
            5'd14:data<=20'b00000000001111100000;
            5'd15:data<=20'b00000000001111000000;
            5'd16:data<=20'b00000000011111000000;
            5'd17:data<=20'b00000000011111000000;
            5'd18:data<=20'b00000000111110000000;
            5'd19:data<=20'b00000000111110000000;
            5'd20:data<=20'b00000000111110000000;
            5'd21:data<=20'b00000001111100000000;
            5'd22:data<=20'b00000001111100000000;
            5'd23:data<=20'b00000011111100000000;
            5'd24:data<=20'b00000011111000000000;
            5'd25:data<=20'b00000011111000000000;
            5'd26:data<=20'b00000111110000000000;
            5'd27:data<=20'b00000111110000000000;
            5'd28:data<=20'b00000111110000000000;
            5'd29:data<=20'b00000111100000000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd8:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000001000000000;
            5'd03:data<=20'b00000011111111000000;
            5'd04:data<=20'b00000111111111100000;
            5'd05:data<=20'b00001111111111110000;
            5'd06:data<=20'b00011111101111111000;
            5'd07:data<=20'b00011111000011111000;
            5'd08:data<=20'b00011110000001111000;
            5'd09:data<=20'b00011110000001111000;
            5'd10:data<=20'b00011110000001111000;
            5'd11:data<=20'b00011111000011111000;
            5'd12:data<=20'b00011111000111110000;
            5'd13:data<=20'b00001111111111100000;
            5'd14:data<=20'b00001111111111100000;
            5'd15:data<=20'b00000111111111000000;
            5'd16:data<=20'b00000011111111000000;
            5'd17:data<=20'b00000111111111110000;
            5'd18:data<=20'b00001111101111110000;
            5'd19:data<=20'b00011111000111111000;
            5'd20:data<=20'b00011110000011111000;
            5'd21:data<=20'b00111110000001111100;
            5'd22:data<=20'b00111100000001111100;
            5'd23:data<=20'b00111100000001111100;
            5'd24:data<=20'b00111110000001111000;
            5'd25:data<=20'b00111111000011111000;
            5'd26:data<=20'b00011111111111111000;
            5'd27:data<=20'b00011111111111110000;
            5'd28:data<=20'b00001111111111100000;
            5'd29:data<=20'b00000011111111000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd9:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000011000000000;
            5'd03:data<=20'b00000011111111000000;
            5'd04:data<=20'b00000111111111100000;
            5'd05:data<=20'b00001111111111110000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011111000011111000;
            5'd08:data<=20'b00111110000011111000;
            5'd09:data<=20'b00111110000001111000;
            5'd10:data<=20'b00111100000001111000;
            5'd11:data<=20'b00111100000001111000;
            5'd12:data<=20'b00111110000001111000;
            5'd13:data<=20'b00111110000001111000;
            5'd14:data<=20'b00111110000001111000;
            5'd15:data<=20'b00011111000111111000;
            5'd16:data<=20'b00011111111111111000;
            5'd17:data<=20'b00011111111111111000;
            5'd18:data<=20'b00001111111111111000;
            5'd19:data<=20'b00000011111001111000;
            5'd20:data<=20'b00000000000001111000;
            5'd21:data<=20'b00000000000001111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011110000;
            5'd24:data<=20'b00000000000111110000;
            5'd25:data<=20'b00011000001111100000;
            5'd26:data<=20'b00011111111111100000;
            5'd27:data<=20'b00011111111111000000;
            5'd28:data<=20'b00011111111110000000;
            5'd29:data<=20'b00001111111000000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd10:
    begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000000000000000;
        5'd04:data<=20'b00000000000000000000;
        5'd05:data<=20'b00000000000000000000;
        5'd06:data<=20'b00000000000000000000;
        5'd07:data<=20'b00000000000000000000;
        5'd08:data<=20'b00000000000000000000;
        5'd09:data<=20'b00000000000000000000;
        5'd10:data<=20'b00000000011111000000;
        5'd11:data<=20'b00000000011111000000;
        5'd12:data<=20'b00000000011111000000;
        5'd13:data<=20'b00000000011111000000;
        5'd14:data<=20'b00000000000000000000;
        5'd15:data<=20'b00000000000000000000;
        5'd16:data<=20'b00000000000000000000;
        5'd17:data<=20'b00000000000000000000;
        5'd18:data<=20'b00000000000000000000;
        5'd19:data<=20'b00000000000000000000;
        5'd20:data<=20'b00000000000000000000;
        5'd21:data<=20'b00000000000000000000;
        5'd22:data<=20'b00000000000000000000;
        5'd23:data<=20'b00000000011111000000;
        5'd24:data<=20'b00000000011111000000;
        5'd25:data<=20'b00000000011111000000;
        5'd26:data<=20'b00000000011111000000;
        5'd27:data<=20'b00000000000000000000;
        5'd28:data<=20'b00000000000000000000;
        5'd29:data<=20'b00000000000000000000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
    end
    default:
        data<=0;    
    endcase
end
always @(posedge clk_25MHz)
begin
    case(data_adrs)
        5'd00:score_t<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd01:score_t<=100'b0000000110000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000;
        5'd02:score_t<=100'b0000111111110000000000011111110000000000011111111100000000001111111110000000001111111111110000000000;
        5'd03:score_t<=100'b0001111111111000000001111111111100000000111111111110000000001111111111100000001111111111110000000000;
        5'd04:score_t<=100'b0011111111111000000011111111111110000001111111111111000000001111111111110000001111111111110000000000;
        5'd05:score_t<=100'b0011100000011000000011110000011110000011110000001111100000001110000011110000001111000000000000000000;
        5'd06:score_t<=100'b0111100000000000000111100000000110000111100000000011100000001110000001111000001110000000000000000000;
        5'd07:score_t<=100'b0111000000000000000111000000000000000111000000000011110000001110000001111000001110000000000000000000;
        5'd08:score_t<=100'b0111000000000000001111000000000000000111000000000001110000001110000000111000001110000000000000000000;
        5'd09:score_t<=100'b0111000000000000001110000000000000001111000000000001110000001110000000111000001110000000000000000000;
        5'd10:score_t<=100'b0111100000000000001110000000000000001110000000000001111000001110000000111000001110000000000000001100;
        5'd11:score_t<=100'b0111100000000000011110000000000000001110000000000000111000001110000000111000001110000000000000001110;
        5'd12:score_t<=100'b0011110000000000011100000000000000001110000000000000111000001110000001111000001110000000000000001110;
        5'd13:score_t<=100'b0011111000000000011100000000000000001110000000000000111000001110000001110000001110000000000000001110;
        5'd14:score_t<=100'b0001111110000000011100000000000000001110000000000000111000001110000111100000001111111111100000001110;
        5'd15:score_t<=100'b0000111111000000011100000000000000001110000000000000111000001111111111100000001111111111100000000000;
        5'd16:score_t<=100'b0000011111110000011100000000000000011110000000000000111000001111111110000000001111111111100000000000;
        5'd17:score_t<=100'b0000000111111000011100000000000000001110000000000000111000001111111111000000001111000000000000000000;
        5'd18:score_t<=100'b0000000011111000011100000000000000001110000000000000111000001110000111000000001110000000000000000000;
        5'd19:score_t<=100'b0000000000111100011100000000000000001110000000000000111000001110000011100000001110000000000000000000;
        5'd20:score_t<=100'b0000000000111100011100000000000000001110000000000000111000001110000011100000001110000000000000000000;
        5'd21:score_t<=100'b0000000000011100011110000000000000001110000000000001111000001110000001110000001110000000000000000000;
        5'd22:score_t<=100'b0000000000011100001110000000000000001110000000000001110000001110000001110000001110000000000000000000;
        5'd23:score_t<=100'b0000000000011100001110000000000000001111000000000001110000001110000001110000001110000000000000000000;
        5'd24:score_t<=100'b0000000000011100001111000000000000000111000000000011110000001110000001111000001110000000000000000000;
        5'd25:score_t<=100'b0000000000011100000111000000000010000111100000000011100000001110000000111000001110000000000000000000;
        5'd26:score_t<=100'b0110000000111000000111100000001110000111100000000111100000001110000000111000001110000000000000001110;
        5'd27:score_t<=100'b0111100001111000000011111000111110000011111000011111000000001110000000111100001111000000000000001110;
        5'd28:score_t<=100'b0111111111110000000011111111111100000001111111111110000000001110000000011100001111111111111000001110;
        5'd29:score_t<=100'b0011111111100000000001111111111000000000111111111100000000001110000000011100001111111111111000001110;
        5'd30:score_t<=100'b0001111111000000000000011111100000000000001111111000000000001110000000011100000111111111111000001110;
        5'd31:score_t<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
end
endmodule

module DATA_DG(clk,data_adrs,data,go_adrs,game_over);
input clk;
input [5:0] data_adrs,go_adrs;
output reg [0:39] data;
output reg [0:235] game_over;
always @(posedge clk)
begin
    case(data_adrs)
        6'd00:data<=40'b0000000000000000000000000000000000000000;
        6'd01:data<=40'b0000000000000000011111111000000000000000;
        6'd02:data<=40'b0000000000000001110011111100000000000000;
        6'd03:data<=40'b0000000000000011001111001100000000000000;
        6'd04:data<=40'b0000000000000001111111111000000000000000;
        6'd05:data<=40'b0000000000000000011111000000000000000000;
        6'd06:data<=40'b0000000000000000000111000000000000000000;
        6'd07:data<=40'b0000000000000000001111100000000000000000;
        6'd08:data<=40'b0000000000000001111111111110000000000000;
        6'd09:data<=40'b0000000000000111111111111111110000000000;
        6'd10:data<=40'b0000000000011111111111111111111000000000;
        6'd11:data<=40'b0000000000111111111100011100011100000000;
        6'd12:data<=40'b0000000001111111111000001000011110000000;
        6'd13:data<=40'b0000000001111111111000001000011111000000;
        6'd14:data<=40'b0000000011111111111001101110011111000000;
        6'd15:data<=40'b0000000011111111111101111110011111100000;
        6'd16:data<=40'b0000000011111111111111111111110111100000;
        6'd17:data<=40'b0000000111111100111111011111111111100000;
        6'd18:data<=40'b0000000111111001111100001110111111100000;
        6'd19:data<=40'b0000000111110001111100001100111111100000;
        6'd20:data<=40'b0000000111110001111111111100111111100000;
        6'd21:data<=40'b0001111111110011111111111111110011100000;
        6'd22:data<=40'b0011001111110011111111111111111110100000;
        6'd23:data<=40'b0010000111110011111111111111111001100000;
        6'd24:data<=40'b0010000111110001111111111111111001000000;
        6'd25:data<=40'b0011001111110000111111111111110011011100;
        6'd26:data<=40'b0001111111110000011111111111100010111110;
        6'd27:data<=40'b0000111111111000001111111111000111100011;
        6'd28:data<=40'b0000111111111000000111111110001111100011;
        6'd29:data<=40'b0000011111111110000001111100011111100010;
        6'd30:data<=40'b0000011111111111111000000111111111111110;
        6'd31:data<=40'b0000001111111111111111111111111111110000;
        6'd32:data<=40'b0000001111111111111111111111111111100000;
        6'd33:data<=40'b0000011111111100000011111001111111000000;
        6'd34:data<=40'b0000011111111000000011111001111110000000;
        6'd35:data<=40'b0000011111110000000001110001111100000000;
        6'd36:data<=40'b0001111111110011111110111111110000000000;
        6'd37:data<=40'b0011011111110010011111111111000000000000;
        6'd38:data<=40'b0010011111110010000000000111000000000000;
        6'd39:data<=40'b0010011111110011000000001110000000000000;
        6'd40:data<=40'b0110011111111001100000111100000000000000;
        6'd41:data<=40'b0110011111111100111111111000000000000000;
        6'd42:data<=40'b0100001111111111111111110000000000000000;
        6'd43:data<=40'b0110000011111111111111100000000000000000;
        6'd44:data<=40'b0010000001011111111110000000000000000000;
        6'd45:data<=40'b0011000111011011111110000000000000000000;
        6'd46:data<=40'b0001111100011000000110000000000000000000;
        6'd47:data<=40'b0000000000001100000100000000000000000000;
        6'd48:data<=40'b0000000000000111111000000000000000000000;
        6'd49:data<=40'b0000000000000001110000000000000000000000;
    endcase
end
always @(posedge clk)
begin
    case(go_adrs)
        6'd00:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd01:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd02:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd03:game_over<=236'b00000000011111111111100000000000000000001111000000000000001111110000000000000000111110000001111111111111111111100000000000000000000000011111111110000000000111100000000000000000011110001111111111111111111100000011111111111111111100000000;
6'd04:game_over<=236'b00000001111111111111111000000000000000011111100000000000001111110000000000000001111110000001111111111111111111100000000000000000000001111111111111100000000011110000000000000000111100001111111111111111111100000011111111111111111111000000;
6'd05:game_over<=236'b00000011111111111111111100000000000000011111100000000000001111111000000000000001111110000001111111111111111111100000000000000000000111111111111111111000000011110000000000000000111100001111111111111111111100000011111111111111111111100000;
6'd06:game_over<=236'b00000111111000000001111110000000000000011111100000000000001111111000000000000001111110000001111000000000000000000000000000000000001111110000000011111100000001111000000000000000111000001111000000000000000000000011110000000000001111100000;
6'd07:game_over<=236'b00001111100000000000011110000000000000111111110000000000001111111000000000000011111110000001111000000000000000000000000000000000011111000000000000111100000001111000000000000001111000001111000000000000000000000011110000000000000111110000;
6'd08:game_over<=236'b00011111000000000000001111000000000000111001110000000000001111111100000000000011111110000001111000000000000000000000000000000000011110000000000000011110000001111000000000000001111000001111000000000000000000000011110000000000000011110000;
6'd09:game_over<=236'b00011110000000000000001111000000000000111001111000000000001111111100000000000011111110000001111000000000000000000000000000000000111100000000000000011111000000111100000000000001110000001111000000000000000000000011110000000000000001110000;
6'd10:game_over<=236'b00111100000000000000000111000000000001111001111000000000001111011100000000000111011110000001111000000000000000000000000000000000111100000000000000001111000000111100000000000011110000001111000000000000000000000011110000000000000001110000;
6'd11:game_over<=236'b00111100000000000000000100000000000001110000111100000000001111011110000000000111011110000001111000000000000000000000000000000001111000000000000000000111000000011100000000000011100000001111000000000000000000000011110000000000000001110000;
6'd12:game_over<=236'b00111100000000000000000000000000000011110000111100000000001111001110000000000111011110000001111000000000000000000000000000000001111000000000000000000111100000011110000000000111100000001111000000000000000000000011110000000000000011110000;
6'd13:game_over<=236'b01111000000000000000000000000000000011110000011100000000001111001110000000001110011110000001111000000000000000000000000000000001111000000000000000000111100000011110000000000111100000001111000000000000000000000011110000000000000011110000;
6'd14:game_over<=236'b01111000000000000000000000000000000011100000011110000000001111001111000000001110011110000001111000000000000000000000000000000001111000000000000000000111100000001110000000000111000000001111000000000000000000000011110000000000001111100000;
6'd15:game_over<=236'b01111000000000000000000000000000000111100000011110000000001111000111000000001110011110000001111111111111111111000000000000000001111000000000000000000111100000001111000000001111000000001111111111111111111000000011111111111111111111100000;
6'd16:game_over<=236'b01111000000000000000000000000000000111000000001111000000001111000111000000011100011110000001111111111111111111000000000000000001110000000000000000000111100000001111000000001111000000001111111111111111111000000011111111111111111110000000;
6'd17:game_over<=236'b01111000000000011111111111100000001111000000001111000000001111000111100000011100011110000001111111111111111111000000000000000001110000000000000000000111100000000111000000001110000000001111111111111111111000000011111111111111111000000000;
6'd18:game_over<=236'b01111000000000011111111111100000001111000000001111000000001111000011100000011100011110000001111000000000000000000000000000000001111000000000000000000111100000000111100000011110000000001111000000000000000000000011111111111111110000000000;
6'd19:game_over<=236'b01111000000000011111111111100000001111111111111111100000001111000011100000111000011110000001111000000000000000000000000000000001111000000000000000000111100000000011100000011100000000001111000000000000000000000011110000000011111000000000;
6'd20:game_over<=236'b01111000000000000000000111100000011111111111111111100000001111000011110000111000011110000001111000000000000000000000000000000001111000000000000000000111100000000011110000011100000000001111000000000000000000000011110000000001111100000000;
6'd21:game_over<=236'b00111100000000000000000111100000011111111111111111110000001111000001110000111000011110000001111000000000000000000000000000000001111000000000000000000111100000000011110000111100000000001111000000000000000000000011110000000000111110000000;
6'd22:game_over<=236'b00111100000000000000000111100000011110000000000011110000001111000001110001110000011110000001111000000000000000000000000000000000111000000000000000000111000000000001110000111000000000001111000000000000000000000011110000000000011110000000;
6'd23:game_over<=236'b00111100000000000000000111100000111100000000000011110000001111000001111001110000011110000001111000000000000000000000000000000000111100000000000000001111000000000001111001111000000000001111000000000000000000000011110000000000011111000000;
6'd24:game_over<=236'b00011110000000000000000111100000111100000000000001111000001111000000111001110000011110000001111000000000000000000000000000000000111110000000000000011111000000000000111001110000000000001111000000000000000000000011110000000000001111100000;
6'd25:game_over<=236'b00011111000000000000000111100001111000000000000001111000001111000000111011100000011110000001111000000000000000000000000000000000011110000000000000011110000000000000111001110000000000001111000000000000000000000011110000000000000111100000;
6'd26:game_over<=236'b00001111100000000000011111100001111000000000000000111100001111000000111111100000011110000001111000000000000000000000000000000000001111100000000001111100000000000000111111110000000000001111000000000000000000000011110000000000000111110000;
6'd27:game_over<=236'b00000111111100000001111111000001110000000000000000111100001111000000011111000000011110000001111000000000000000000000000000000000000111110000000011111100000000000000011111100000000000001111000000000000000000000011110000000000000011111000;
6'd28:game_over<=236'b00000011111111111111111110000011110000000000000000111110001111000000011111000000011110000001111111111111111111110000000000000000000011111111111111110000000000000000011111100000000000001111111111111111111110000011110000000000000001111000;
6'd29:game_over<=236'b00000000111111111111111000000011110000000000000000011110001111000000011111000000011110000001111111111111111111110000000000000000000001111111111111100000000000000000001111000000000000001111111111111111111110000011110000000000000001111100;
6'd30:game_over<=236'b00000000001111111111100000000011100000000000000000011110001111000000001110000000011110000001111111111111111111110000000000000000000000011111111110000000000000000000001111000000000000001111111111111111111110000011110000000000000000111100;
6'd31:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd32:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd33:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd34:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd35:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd36:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd37:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd38:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd39:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd40:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd41:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd42:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd43:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110111000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd44:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110111000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd45:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd46:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd47:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd48:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd49:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd50:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd51:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd52:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd53:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd54:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd55:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd56:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd57:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd58:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd59:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd60:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd61:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd62:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd63:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
end
endmodule