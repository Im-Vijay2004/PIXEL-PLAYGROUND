module DODGE_CAR(sys_clk,clk_25M,rt,lt,reset1,hcount,vcount,red,green,blue,rst_dc);
input sys_clk,clk_25M;
input rt,lt,reset1,rst_dc;
input[9:0] hcount,vcount;
output [3:0] red,green,blue;
wire [9:0] hcount,vcount;
wire clk_100,clk_50,clk_10,clk_02,stop;

wire [5:0] data_adrs,go_adrs,tree_adrs1,obs_adrs1,tree_adrs2,obs_adrs2,tree_adrs3,obs_adrs3,tree_adrs4,obs_adrs4,tree_adrs5,obs_adrs5,tree_adrs6,obs_adrs6,tree_adrs7,obs_adrs7;
wire [4:0] score_adrs;
wire [0:235] game_over;
wire [0:31] data,obstacle1,obstacle2,obstacle3,obstacle4,obstacle5,obstacle6,obstacle7;
wire [0:49] tree1,tree2,tree3,tree4,tree5,tree6;
wire stop_temp;
wire [0:19] score1,score2,score3,score4;
wire [3:0] bcd3,bcd2,bcd1,bcd0;
wire [15:0] bcd;
wire [0:99] score_t;
assign bcd3=bcd[15:12];
assign bcd2=bcd[11:8];
assign bcd1=bcd[7:4];
assign bcd0=bcd[3:0];
assign stop_temp=0;
wire reset;
assign reset=reset1|rst_dc;
CLK_100Hz_DC clk_div2(sys_clk,clk_100);
CLK_02Hz_DC clk_div3(sys_clk,clk_02);
CLK_10Hz_DC clk_div4(sys_clk,clk_10);
CLK_50Hz_DC clk_div5(sys_clk,clk_50);
DISP_WRITE_DC disp(clk_25M,clk_100,clk_50,clk_02,hcount,vcount,red,green,blue,rt,lt,reset,score1,score2,score3,score4,score_t,score_adrs,stop,data_adrs,data,score_adrs,go_adrs,game_over,tree_adrs1,tree_adrs2,tree_adrs3,tree_adrs4,tree_adrs5,tree_adrs6,tree1,tree2,tree3,tree4,tree5,tree6,obs_adrs1,obs_adrs2,obs_adrs3,obs_adrs4,obs_adrs5,obs_adrs6,obs_adrs7,obstacle1,obstacle2,obstacle3,obstacle4,obstacle5,obstacle6,obstacle7);
SCORE_DC Score_counter(sys_clk,bcd,stop,reset);
SCORE_DATA_DC Score1(clk_25M,bcd0,score1,score_adrs,score_t);
SCORE_DATA_DC Score2(clk_25M,bcd1,score2,score_adrs);
SCORE_DATA_DC Score3(clk_25M,bcd2,score3,score_adrs);
SCORE_DATA_DC Score4(clk_25M,bcd3,score4,score_adrs);


MAIN_DATA_DC Car(clk_25M,data_adrs,data,go_adrs,game_over);
TREE_OBSTACLE_DC TOBS(clk_25M,obs_adrs1,obstacle1,tree_adrs1,tree1);
TREE_OBSTACLE_DC TOBS2(clk_25M,obs_adrs2,obstacle2,tree_adrs2,tree2);
TREE_OBSTACLE_DC TOBS3(clk_25M,obs_adrs3,obstacle3,tree_adrs3,tree3);
TREE_OBSTACLE_DC TOBS4(clk_25M,obs_adrs4,obstacle4,tree_adrs4,tree4);
TREE_OBSTACLE_DC TOBS5(clk_25M,obs_adrs5,obstacle5,tree_adrs5,tree5);
TREE_OBSTACLE_DC TOBS6(clk_25M,obs_adrs6,obstacle6,tree_adrs6,tree6);
TREE_OBSTACLE_DC TOBS7(clk_25M,obs_adrs7,obstacle7,tree_adrs7,tree7);

endmodule

module CLK_100Hz_DC(clk_in,clk_out);
input clk_in;
output reg clk_out=0;
integer i;
always @(posedge clk_in)
begin
    if(i==499999)
    begin
        clk_out<=~clk_out;
        i<=0;
    end
    else
        i<=i+1;
end
endmodule


module CLK_02Hz_DC(clk_in,clk_out);
input clk_in;
output reg clk_out=0;
integer i;
always @(posedge clk_in)
begin
    if(i==249999999)
    begin
        clk_out<=~clk_out;
        i<=0;
    end
    else
        i<=i+1;
end
endmodule
module CLK_10Hz_DC(clk_in,clk_out);
input clk_in;
output reg clk_out=0;
integer i;
always @(posedge clk_in)
begin
    if(i==4999999)
    begin
        clk_out<=~clk_out;
        i<=0;
    end
    else
        i<=i+1;
end
endmodule
module CLK_50Hz_DC(clk_in,clk_out);
input clk_in;
output reg clk_out=0;
integer i;
always @(posedge clk_in)
begin
    if(i==999998)
    begin
        clk_out<=~clk_out;
        i<=0;
    end
    else
        i<=i+1;
end
endmodule

module DISP_WRITE_DC(clk_25M,clk_100,clk_50,clk_02,hcount,vcount,red,green,blue,push_right,push_left,rst,score1,score2,score3,score4,score_t,score_adrs,stop,data_adrs,data,score_adrs,go_adrs,game_over,tree_adrs1,tree_adrs2,tree_adrs3,tree_adrs4,tree_adrs5,tree_adrs6,tree1,tree2,tree3,tree4,tree5,tree6,obs_adrs1,obs_adrs2,obs_adrs3,obs_adrs4,obs_adrs5,obs_adrs6,obs_adrs7,obstacle1,obstacle2,obstacle3,obstacle4,obstacle5,obstacle6,obstacle7);
input clk_25M,push_right,push_left,clk_100,clk_50,clk_02,rst;
input [0:19] score1;
input [0:19] score2;
input [0:19] score3;
input [0:19] score4;
input [0:99] score_t;
output reg stop;
input [0:31] data,obstacle1,obstacle2,obstacle3,obstacle4,obstacle5,obstacle6,obstacle7;
input [0:49] tree1;
input [0:49] tree2;
input [0:49] tree3;
input [0:49] tree4;
input [0:49] tree5;
input [0:49] tree6;
output reg [5:0] data_adrs,obs_adrs1,obs_adrs2,obs_adrs3,obs_adrs4,obs_adrs5,obs_adrs6,obs_adrs7;
output reg [5:0] go_adrs;
output reg [5:0] tree_adrs1;
output reg [5:0] tree_adrs2;
output reg [5:0] tree_adrs3;
output reg [5:0] tree_adrs4;
output reg [5:0] tree_adrs5;
output reg [5:0] tree_adrs6;
output reg [4:0] score_adrs;
input [0:235] game_over;
input [9:0] hcount,vcount;

reg [9:0]move=275;
reg [9:0]temp=514;
reg [9:0]up1=0;
reg [9:0]up2=65;
reg [9:0]up3=130;
reg [9:0]up4=195;
reg [9:0]up5=260;
reg [9:0]up6=325;
reg [9:0]up7=390;
reg [9:0]up8=455;
reg [8:0]tree_move1=85;
reg [8:0]tree_move2=245;
reg [8:0]tree_move3=405;
reg [8:0]tree_move4=85;
reg [8:0]tree_move5=245;
reg [8:0]tree_move6=405;


output reg [3:0] red,green,blue;
parameter   hmin=144,
            hmax=784,
            vmin=35,
            vmax=515,
            box1=314,
            box2=465;            
            reg [9:0]obs1=0;
            reg [9:0]obs2=150;
            reg [9:0]obs3=300;
            reg [9:0]obs4=450;
            reg [9:0]obs5=600;
            reg [9:0]obs6=750;
            reg [9:0]obs7=900;
            
always @(posedge clk_25M)
begin
    if((hcount>=hmin && hcount<=hmax) && (vcount>=vmin && vcount<=vmax))
        begin
        data_adrs<=vcount-move;
        //data_adrs<=hcount-temp;
         score_adrs<=vcount-40;
          go_adrs<=vcount-263;
          tree_adrs1<=vcount-tree_move1;
           tree_adrs2<=vcount-tree_move2;
            tree_adrs3<=vcount-tree_move3;
             tree_adrs4<=vcount-tree_move4;
              tree_adrs5<=vcount-tree_move5;
               tree_adrs6<=vcount-tree_move6;
               obs_adrs1<=vcount-obs1;
               obs_adrs2<=vcount-obs2;
               obs_adrs3<=vcount-obs3;
               obs_adrs4<=vcount-obs4;
               obs_adrs5<=vcount-obs5;
               obs_adrs6<=vcount-obs6;
               obs_adrs7<=vcount-obs7;
               
                 if((hcount>=346 && hcount<=582) && (vcount>=263 && vcount<=327)&&(game_over[hcount-346]==1)&& stop)//gameover
            begin
                {red,green,blue}<={4'b1111,4'b0000,4'b0000};
            end
         else if((hcount>=temp && hcount<=temp+32) && (vcount>=move && vcount<=move+50) && (data[hcount-temp]==1))//car
                begin
                     {red,green,blue}<={4'b1111,4'b0000,4'b0000};
                end
           else if((hcount>=750 && hcount<=770) && (vcount>=40 && vcount<=72)&&(score1[hcount-750]==1))
            begin
                {red,green,blue}<={4'b1100,4'b1110,4'b1110};
            end
            else if((hcount>=730 && hcount<=750) && (vcount>=40 && vcount<=72)&&(score2[hcount-730]==1))
            begin
                {red,green,blue}<={4'b1100,4'b1110,4'b1110};
            end
            else if((hcount>=710 && hcount<=730) && (vcount>=40 && vcount<=72) && (score3[hcount-710]==1))
            begin
                {red,green,blue}<={4'b1100,4'b1110,4'b1110};
            end
            else if((hcount>=690 && hcount<=710) && (vcount>=40 && vcount<=72)&&(score4[hcount-690]==1))
            begin
                {red,green,blue}<={4'b1100,4'b1110,4'b1110};
            end
            else if((hcount>=590 && hcount<=689) && (vcount>=40 && vcount<=72)&&(score_t[hcount-590]==1))
            begin
                {red,green,blue}<={4'b1100,4'b1110,4'b1110};
            end
            else if((hcount>=150 && hcount<=200) && (vcount>=tree_move1 && vcount<=tree_move1+60) && (tree1[hcount-150]==1))//left_tree-1
                begin
                     {red,green,blue}<={4'b0000,4'b1111,4'b0000};
                end
            else if((hcount>=240 && hcount<=290) && (vcount>=tree_move2 && vcount<=tree_move2+60)&& (tree2[hcount-240]==1))//left_tree-2
                begin
                     {red,green,blue}<={4'b0000,4'b1111,4'b0000};
                end
             else if((hcount>=150 && hcount<=200) && (vcount>=tree_move3 && vcount<=tree_move3+60) && (tree3[hcount-150]==1))//left_tree-3
                begin
                     {red,green,blue}<={4'b0000,4'b1111,4'b0000};
                end
             else if((hcount>=720 && hcount<=770) && (vcount>=tree_move4 && vcount<=tree_move4+60) && (tree4[hcount-720]==1))//right_tree-1
                begin
                     {red,green,blue}<={4'b0000,4'b1111,4'b0000};
                end
            else if((hcount>=630 && hcount<=680) && (vcount>=tree_move5 && vcount<=tree_move5+60)&& (tree5[hcount-630]==1))//right_tree-2
                begin
                     {red,green,blue}<={4'b0000,4'b1111,4'b0000};
                end
                 else if((hcount>=720 && hcount<=770) && (vcount>=tree_move6 && vcount<=tree_move6+60) && (tree6[hcount-720]==1))//right tree-3
            begin
                {red,green,blue}<={4'b0000,4'b1111,4'b0000};
            end
          else if((hcount>=364 && hcount<=396) && (vcount>=obs1 && vcount<=obs1+50) && (obstacle1[hcount-364]==1))//obstacle-1
                begin
                     {red,green,blue}<={4'b0000,4'b0000,4'b1111};
                end
          else if((hcount>=514 && hcount<=546) && (vcount>=obs2 && vcount<=obs2+50) && (obstacle2[hcount-514]==1))//obstacle-2
                begin
                     {red,green,blue}<={4'b1111,4'b1100,4'b1110};
                end
                 else if((hcount>=364 && hcount<=396) && (vcount>=obs3 && vcount<=obs3+50)&& (obstacle3[hcount-364]==1))//obstacle-3
                begin
                     {red,green,blue}<={4'b1110,4'b1110,4'b0100};
                end
          else if((hcount>=514 && hcount<=546) && (vcount>=obs4 && vcount<=obs4+50)&& (obstacle4[hcount-514]==1) )//obstacle-4
                begin
                     {red,green,blue}<={4'b0000,4'b0000,4'b1111};
                end
             else if((hcount>=364 && hcount<=396) && (vcount>=obs5 && vcount<=obs5+50) && (obstacle5[hcount-364]==1))//obstacle-5
                begin
                     {red,green,blue}<={4'b1111,4'b1100,4'b1110};
                end
             else if((hcount>=514 && hcount<=546) && (vcount>=obs6 && vcount<=obs6+50) && (obstacle6[hcount-514]==1))//obstacle-6
                begin
                     {red,green,blue}<={4'b1110,4'b1110,4'b0100};
                end
             else if((hcount>=364 && hcount<=396) && (vcount>=obs7 && vcount<=obs7+50) && (obstacle7[hcount-364]==1))//obstacle-7
                begin
                     {red,green,blue}<={4'b0000,4'b0000,4'b1111};
                end
            else if((hcount>=461 && hcount<=467) && (vcount>=up1 && vcount<=up1+65))// first line
                begin
                     {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                end
          else if((hcount>=461 && hcount<=467) && (vcount>=up2 && vcount<=up2+65))//secnd-line-white
                begin
                     {red,green,blue}<={4'b0000,4'b0000,4'b0000};
                end
           else if((hcount>=461 && hcount<=467) && (vcount>=up3 && vcount<=up3+65))//3rd line-black
                begin
                     {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                end
            else if((hcount>=461 && hcount<=467) && (vcount>=up4 && vcount<=up4+65))//4thline-white
                begin
                     {red,green,blue}<={4'b0000,4'b0000,4'b0000};
                end  
             else if((hcount>=461 && hcount<=467) && (vcount>=up5 && vcount<=up5+65))//5th line-black
                begin
                     {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                end  
             else if((hcount>=461 && hcount<=467) && (vcount>=up6 && vcount<=up6+65))//6th line-black
                begin
                     {red,green,blue}<={4'b0000,4'b0000,4'b0000};
                end  
             else if((hcount>=461 && hcount<=467) && (vcount>=up7 && vcount<=up7+65))//7th line-black
                begin
                     {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                end 
             else if((hcount>=461 && hcount<=467) && (vcount>=up8 && vcount<=up8+65))//8th line-black
                begin
                     {red,green,blue}<={4'b0000,4'b0000,4'b0000};
                end   
             else if((hcount>=hmin && hcount<=hmin+170) && (vcount>=35 && vcount<=521))
                begin
                    {red,green,blue}<={4'b1001,4'b1010,4'b1010};
                end
           
            else if((hcount>614 && hcount<=784) && (vcount>=35 && vcount<=521))
                begin
                    {red,green,blue}<={4'b1001,4'b1010,4'b1010};
                end
            else 
                begin
                    {red,green,blue}<={4'b0000,4'b0000,4'b0000};
                end
            end
         else
            begin
                {red,green,blue}<={4'b0000,4'b0000,4'b0000};
            end            
end
//--------------------------CAR movement-----------------------
always@(posedge clk_100)
begin
    if(rst)
        temp<=514;
    else if(!stop)
    begin
    if(temp<box2 && temp>box1)
    begin
        if(push_right)
            temp<=514;
       else if(push_left)
            temp<=temp;
        else
            temp<=temp;
    end
     if(temp<614 && temp>box2)
    begin
        if(push_right)
            temp<=temp;
        else if(push_left)
             temp<=364;
        else
            temp<=temp;
    end
end
end
//--------------------------------white lines movemnet-----------------------
always@(posedge clk_100)
begin
if(!stop && !rst)
begin
     if(up1>515)
        up1<=0;
     else if(up2>515)
        up2<=0;
    else if(up3>515)
        up3<=0;
    else if(up4>515)
        up4<=0;
    else if(up5>515)
        up5<=0;
    else if(up6>515)
        up6<=0;
    else if(up7>515)
        up7<=0;
     else if(up8>515)
        up8<=0;
     else
        begin
            up1<=up1+1;
            up2<=up2+1;
            up3<=up3+1;
            up4<=up4+1;
            up5<=up5+1;
            up6<=up6+1;
            up7<=up7+1;
            up8<=up8+1;
      end 
end
end
//---------------------------stop logic---------------------------
always@(posedge clk_100)
 begin
    if(((temp>=364 && temp <=396) && ((move>=obs1 && move<=obs1+50) || (move+50>=obs1 && move+50<=obs1+50)))||  
    ((temp>=364 && temp <=396) && ((move>=obs3 && move<=obs3+50) || (move+50>=obs3 && move+50<=obs3+50)))||  
    ((temp>=364 && temp <=396) && ((move>=obs5 && move<=obs5+50) || (move+50>=obs5 && move+50<=obs5+50)))|| 
    ((temp>=364 && temp <=396) && ((move>=obs7 && move<=obs7+50) || (move+50>=obs7 && move+50<=obs7+50)))||  
    ((temp>=514 && temp<=546) && ((move>=obs2 && move<=obs2+50) || (move+50>=obs2 && move+50<=obs2+50))) ||  
    ((temp>=514 && temp<=546) && ((move>=obs4 && move<=obs4+50) || (move+50>=obs4 && move+50<=obs4+50))) || 
     ((temp>=514 && temp<=546) && ((move>=obs6 && move<=obs6+50) || (move+50>=obs6 && move+50<=obs6+50))))
     begin
        stop<=1;
        if(rst)
        begin
            stop<=0;
        end
     end
     else
        stop=0;
     end
 //---------------------obstacle movemnet---------------------------
 always@(posedge clk_50)
 begin
 if(!stop)
  begin
        if(rst)
        begin
        obs1<=0; 
        obs2<=150;
        obs3<=300;
        obs4<=450;
        obs5<=600;
        obs6<=750;
        obs7<=900;
        tree_move1<=85; 
        tree_move2<=245;
        tree_move3<=405;
        tree_move4<=85; 
        tree_move5<=245;
        tree_move6<=405;
        end
        else
        begin
        obs1<=obs1+1;
        obs2<=obs2+1;
        obs3<=obs3+1;
        obs4<=obs4+1;
        obs5<=obs5+1;
        obs6<=obs6+1;
        obs7<=obs7+1;
        tree_move1<=tree_move1+1;
        tree_move2<=tree_move2+1;
        tree_move3<=tree_move3+1;
        tree_move4<=tree_move4+1;
        tree_move5<=tree_move5+1;
        tree_move6<=tree_move6+1;
        end
        end
//        else
//        begin
//        if(rst)
//        begin
//        obs1<=0; 
//        obs2<=150;
//        obs3<=300;
//        obs4<=450;
//        obs5<=600;
//        obs6<=750;
//        obs7<=900;
//        tree_move1<=85; 
//        tree_move2<=245;
//        tree_move3<=405;
//        tree_move4<=85; 
//        tree_move5<=245;
//        tree_move6<=405;
//        end
//     else
//        obs1<=obs1; 
//        obs2<=obs2;
//        obs4<=obs4;
//        obs5<=obs5;
//        obs6<=obs6;
//        obs7<=obs7;
//        tree_move1<=tree_move1; 
//        tree_move2<=tree_move2;
//        tree_move3<=tree_move3;
//        tree_move4<=tree_move4; 
//        tree_move5<=tree_move5;
//        tree_move6<=tree_move6;
//        end
end
endmodule


module SCORE_DC(clk,score,stop_temp,reset);
input clk,reset,stop_temp;
output [15:0] score;
reg clk_div;
integer i;
integer div;
reg [13:0] bin=0;
always @(posedge clk)
begin
    if(i==div)
    begin
        clk_div<=~clk_div;
        i<=0;
    end
    else
        i<=i+1;
end
always @(posedge clk)
begin
    if(bin <15)
        div<=49999999;
    else if( bin>=15 && bin <=30)
        div<=25999999;
    else if( bin>30 && bin <=50)
        div<=12599999;
    else if( bin>50 && bin <=100)
        div<=10000000;
    else if( bin>100 && bin <=1000)
        div<=4999999;
    else if( bin>1000 && bin <10000)
        div<=2599999;
    else
        div<=div;
end
always @(posedge clk_div, posedge reset)
begin
    if(reset)
        bin<=0;
    else if(stop_temp)
        bin<=bin;
    else
        bin<=bin+1;
end
BIN_BCD_DC Binary_BCD(clk,bin,score);
endmodule

module BIN_BCD_DC(
input clk,
input [13:0]bin,
output reg [15:0]bcd
);
reg [3:0]count=0;
reg [15:0] bcd_temp=0;
reg reset=0;
always@(posedge clk)
if(reset) begin
    bcd_temp=0;
    count=0;
    reset=0;
end
else if(count<=13)
begin
    if(bcd_temp[3:0]>=5) bcd_temp[3:0]=bcd_temp[3:0]+3;
    if(bcd_temp[7:4]>=5) bcd_temp[7:4]=bcd_temp[7:4]+3;
    if(bcd_temp[11:8]>=5) bcd_temp[11:8]=bcd_temp[11:8]+3;
    if(bcd_temp[15:12]>=5) bcd_temp[15:12]=bcd_temp[15:12]+3;
    bcd_temp={bcd_temp[14:0],bin[13-count]};
    count=count+1;
end
else
begin
    reset=1;
    bcd=bcd_temp;
end
endmodule
module MAIN_DATA_DC(clk,data_adrs,data,go_adrs,game_over);
input clk;
input [5:0] data_adrs,go_adrs;
output reg [0:31] data;
output reg [0:235] game_over;
always @(posedge clk)                                           //car
begin
    case(data_adrs)
        6'd00:data<=32'b0000000000111111111111111100000;
        6'd01:data<=32'b0000000000111111111111111100000;
        6'd02:data<=32'b0000000000111111111111111100000;
        6'd03:data<=32'b0000000000111111111111111100000;
        6'd04:data<=32'b0000000001011111000011111010000;
        6'd05:data<=32'b0000000001111111000011111111000;
        6'd06:data<=32'b0000000001011111000011111011000;
        6'd07:data<=32'b0000000011011111000011111011000;
        6'd08:data<=32'b0000000111011101000010111011100;
        6'd09:data<=32'b0000000111111101000010111011100;
        6'd10:data<=32'b0000000101111101000010111111100;
        6'd11:data<=32'b0000000111111111000011111111100;
        6'd12:data<=32'b0000000111111111000011111111100;
        6'd13:data<=32'b0000000111111111000011111111100;
        6'd14:data<=32'b0000000011111111000011111111100;
        6'd15:data<=32'b0000000011111111111111111111000;
        6'd16:data<=32'b0000000001111000000000011111000;
        6'd17:data<=32'b0000000001110000000000000111000;
        6'd18:data<=32'b0000000001100000000000000111000;
        6'd19:data<=32'b0000000010110000000000000101000;
        6'd20:data<=32'b0000000011111000000000001111100;
        6'd21:data<=32'b0000000011111111111111111111000;
        6'd22:data<=32'b0000000001110111000011111111000;
        6'd23:data<=32'b0000000001111111000011111011000;
        6'd24:data<=32'b0000000001111111000011111011000;
        6'd25:data<=32'b0000000001111111000011111011000;
        6'd26:data<=32'b0000000001111111000011111011000;
        6'd27:data<=32'b0000000001111111000011111111000;
        6'd28:data<=32'b0000000011111111000011111111000;
        6'd29:data<=32'b0000000011111111000011111011000;
        6'd30:data<=32'b0000000001111111000011111011000;
        6'd31:data<=32'b0000000001111111000011111011000;
        6'd32:data<=32'b0000000001111111000011111111000;
        6'd33:data<=32'b0000000011111111000011111111000;
        6'd34:data<=32'b0000000101111111111111111111100;
        6'd35:data<=32'b0000000101111000000110011111100;
        6'd36:data<=32'b0000000101111000001110001111100;
        6'd37:data<=32'b0000000111110000000000001111100;
        6'd38:data<=32'b0000000111110000000000001111100;
        6'd39:data<=32'b0000000111110000000000001111100;
        6'd40:data<=32'b0000000111111111111111111111100;
        6'd41:data<=32'b0000000011111111001011111111000;
        6'd42:data<=32'b0000000001111111111111111111000;
        6'd43:data<=32'b0000000001111111111111111111000;
        6'd44:data<=32'b0000000001111111111111111110000;
        6'd45:data<=32'b0000000001111111111111111110000;
        6'd46:data<=32'b0000000000111111111111111100000;
        6'd47:data<=32'b0000000000111111111111111100000;
        6'd48:data<=32'b0000000000111111111111111100000;
        6'd49:data<=32'b0000000000111111111111111100000;
    endcase
end


always @(posedge clk)
begin
    case(go_adrs)
6'd00:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd01:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd02:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd03:game_over<=236'b00000000011111111111100000000000000000001111000000000000001111110000000000000000111110000001111111111111111111100000000000000000000000011111111110000000000111100000000000000000011110001111111111111111111100000011111111111111111100000000;
6'd04:game_over<=236'b00000001111111111111111000000000000000011111100000000000001111110000000000000001111110000001111111111111111111100000000000000000000001111111111111100000000011110000000000000000111100001111111111111111111100000011111111111111111111000000;
6'd05:game_over<=236'b00000011111111111111111100000000000000011111100000000000001111111000000000000001111110000001111111111111111111100000000000000000000111111111111111111000000011110000000000000000111100001111111111111111111100000011111111111111111111100000;
6'd06:game_over<=236'b00000111111000000001111110000000000000011111100000000000001111111000000000000001111110000001111000000000000000000000000000000000001111110000000011111100000001111000000000000000111000001111000000000000000000000011110000000000001111100000;
6'd07:game_over<=236'b00001111100000000000011110000000000000111111110000000000001111111000000000000011111110000001111000000000000000000000000000000000011111000000000000111100000001111000000000000001111000001111000000000000000000000011110000000000000111110000;
6'd08:game_over<=236'b00011111000000000000001111000000000000111001110000000000001111111100000000000011111110000001111000000000000000000000000000000000011110000000000000011110000001111000000000000001111000001111000000000000000000000011110000000000000011110000;
6'd09:game_over<=236'b00011110000000000000001111000000000000111001111000000000001111111100000000000011111110000001111000000000000000000000000000000000111100000000000000011111000000111100000000000001110000001111000000000000000000000011110000000000000001110000;
6'd10:game_over<=236'b00111100000000000000000111000000000001111001111000000000001111011100000000000111011110000001111000000000000000000000000000000000111100000000000000001111000000111100000000000011110000001111000000000000000000000011110000000000000001110000;
6'd11:game_over<=236'b00111100000000000000000100000000000001110000111100000000001111011110000000000111011110000001111000000000000000000000000000000001111000000000000000000111000000011100000000000011100000001111000000000000000000000011110000000000000001110000;
6'd12:game_over<=236'b00111100000000000000000000000000000011110000111100000000001111001110000000000111011110000001111000000000000000000000000000000001111000000000000000000111100000011110000000000111100000001111000000000000000000000011110000000000000011110000;
6'd13:game_over<=236'b01111000000000000000000000000000000011110000011100000000001111001110000000001110011110000001111000000000000000000000000000000001111000000000000000000111100000011110000000000111100000001111000000000000000000000011110000000000000011110000;
6'd14:game_over<=236'b01111000000000000000000000000000000011100000011110000000001111001111000000001110011110000001111000000000000000000000000000000001111000000000000000000111100000001110000000000111000000001111000000000000000000000011110000000000001111100000;
6'd15:game_over<=236'b01111000000000000000000000000000000111100000011110000000001111000111000000001110011110000001111111111111111111000000000000000001111000000000000000000111100000001111000000001111000000001111111111111111111000000011111111111111111111100000;
6'd16:game_over<=236'b01111000000000000000000000000000000111000000001111000000001111000111000000011100011110000001111111111111111111000000000000000001110000000000000000000111100000001111000000001111000000001111111111111111111000000011111111111111111110000000;
6'd17:game_over<=236'b01111000000000011111111111100000001111000000001111000000001111000111100000011100011110000001111111111111111111000000000000000001110000000000000000000111100000000111000000001110000000001111111111111111111000000011111111111111111000000000;
6'd18:game_over<=236'b01111000000000011111111111100000001111000000001111000000001111000011100000011100011110000001111000000000000000000000000000000001111000000000000000000111100000000111100000011110000000001111000000000000000000000011111111111111110000000000;
6'd19:game_over<=236'b01111000000000011111111111100000001111111111111111100000001111000011100000111000011110000001111000000000000000000000000000000001111000000000000000000111100000000011100000011100000000001111000000000000000000000011110000000011111000000000;
6'd20:game_over<=236'b01111000000000000000000111100000011111111111111111100000001111000011110000111000011110000001111000000000000000000000000000000001111000000000000000000111100000000011110000011100000000001111000000000000000000000011110000000001111100000000;
6'd21:game_over<=236'b00111100000000000000000111100000011111111111111111110000001111000001110000111000011110000001111000000000000000000000000000000001111000000000000000000111100000000011110000111100000000001111000000000000000000000011110000000000111110000000;
6'd22:game_over<=236'b00111100000000000000000111100000011110000000000011110000001111000001110001110000011110000001111000000000000000000000000000000000111000000000000000000111000000000001110000111000000000001111000000000000000000000011110000000000011110000000;
6'd23:game_over<=236'b00111100000000000000000111100000111100000000000011110000001111000001111001110000011110000001111000000000000000000000000000000000111100000000000000001111000000000001111001111000000000001111000000000000000000000011110000000000011111000000;
6'd24:game_over<=236'b00011110000000000000000111100000111100000000000001111000001111000000111001110000011110000001111000000000000000000000000000000000111110000000000000011111000000000000111001110000000000001111000000000000000000000011110000000000001111100000;
6'd25:game_over<=236'b00011111000000000000000111100001111000000000000001111000001111000000111011100000011110000001111000000000000000000000000000000000011110000000000000011110000000000000111001110000000000001111000000000000000000000011110000000000000111100000;
6'd26:game_over<=236'b00001111100000000000011111100001111000000000000000111100001111000000111111100000011110000001111000000000000000000000000000000000001111100000000001111100000000000000111111110000000000001111000000000000000000000011110000000000000111110000;
6'd27:game_over<=236'b00000111111100000001111111000001110000000000000000111100001111000000011111000000011110000001111000000000000000000000000000000000000111110000000011111100000000000000011111100000000000001111000000000000000000000011110000000000000011111000;
6'd28:game_over<=236'b00000011111111111111111110000011110000000000000000111110001111000000011111000000011110000001111111111111111111110000000000000000000011111111111111110000000000000000011111100000000000001111111111111111111110000011110000000000000001111000;
6'd29:game_over<=236'b00000000111111111111111000000011110000000000000000011110001111000000011111000000011110000001111111111111111111110000000000000000000001111111111111100000000000000000001111000000000000001111111111111111111110000011110000000000000001111100;
6'd30:game_over<=236'b00000000001111111111100000000011100000000000000000011110001111000000001110000000011110000001111111111111111111110000000000000000000000011111111110000000000000000000001111000000000000001111111111111111111110000011110000000000000000111100;
6'd31:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd32:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd33:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd34:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd35:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd36:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd37:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd38:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd39:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd40:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd41:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd42:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd43:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110111000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd44:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110111000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd45:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd46:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd47:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd48:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd49:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd50:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd51:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd52:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd53:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd54:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd55:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd56:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd57:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd58:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd59:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd60:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd61:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd62:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd63:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
end
endmodule

module TREE_OBSTACLE_DC(clk,obs_adrs,obs,tree_adrs,tree);
input clk;
input [5:0] obs_adrs,tree_adrs;
output reg [31:0] obs;
output reg [49:0] tree;
always @(posedge clk)
begin
    case(tree_adrs)
        6'd00:tree<=50'b00000000000000000000000000011111100000000000000000;
        6'd01:tree<=50'b00000000000000000000010000011111110000000000000000;
        6'd02:tree<=50'b00000000000000001111111101111111111100000000000000;
        6'd03:tree<=50'b00000000000000111111111111111111111110000000000000;
        6'd04:tree<=50'b00000000000000111111111111111111111111110000000000;
        6'd05:tree<=50'b00000000000111111111111111111111111111110000000000;
        6'd06:tree<=50'b00000000001111111111111111111111111111111000000000;
        6'd07:tree<=50'b00000000011111111111111111111111111111111000000000;
        6'd08:tree<=50'b00000001111111111111111111111111111111111100000000;
        6'd09:tree<=50'b00000001111111111111111111111111111111111100000000;
        6'd10:tree<=50'b00000001111111111111111111111111111111111100000000;
        6'd11:tree<=50'b00000001111111111111111111111111111111111110000000;
        6'd12:tree<=50'b00000001111111111111111111111111111111111111000000;
        6'd13:tree<=50'b00000111111111111111111111111111111111111111100000;
        6'd14:tree<=50'b00000111111111111111111111111111111111111111100000;
        6'd15:tree<=50'b00001111111111111111111111111111111111111111110000;
        6'd16:tree<=50'b00000111111111111111111111111111111111111111111000;
        6'd17:tree<=50'b01111111111111111111111111111111111111111111111100;
        6'd18:tree<=50'b01111111111111111111111111111111111111111111111110;
        6'd19:tree<=50'b11111111111111111111111111111111111111111111111110;
        6'd20:tree<=50'b01111111111111111111111111111111111111111111111110;
        6'd21:tree<=50'b00011111111111111111111111111111111111111111111110;
        6'd22:tree<=50'b00011110111111111111111111111111110111111111111100;
        6'd23:tree<=50'b00000010010011111111110111111111000110111111111100;
        6'd24:tree<=50'b00000000000000011000001111001000000011111111111000;
        6'd25:tree<=50'b00000000000000000000000111010000000011110011000000;
        6'd26:tree<=50'b00000000000000000000000011100000000000000000000000;
        6'd27:tree<=50'b00000000000000000000000011000000000000000000000000;
        6'd28:tree<=50'b00000000000000000000000011000000000000000000000000;
        6'd29:tree<=50'b00000000000000000000000011000000000000000000000000;
        6'd30:tree<=50'b00000000000000000000000011100000000000000000000000;
        6'd31:tree<=50'b00000000000000000000000011100000000000000000000000;
        6'd32:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd33:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd34:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd35:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd36:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd37:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd38:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd39:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd40:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd41:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd42:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd43:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd44:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd45:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd46:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd47:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd48:tree<=50'b00000000000000000000011111111100000000000000000000;
        6'd49:tree<=50'b00000000000000000000011111111100000000000000000000;
    endcase             
end

always @(posedge clk)                                           //car
begin
    case(obs_adrs)
        6'd00:obs<=32'b0000000000111111111111111100000;
        6'd01:obs<=32'b0000000000111111111111111100000;
        6'd02:obs<=32'b0000000000111111111111111100000;
        6'd03:obs<=32'b0000000000111111111111111100000;
        6'd04:obs<=32'b0000000001011111000011111010000;
        6'd05:obs<=32'b0000000001111111000011111111000;
        6'd06:obs<=32'b0000000001011111000011111011000;
        6'd07:obs<=32'b0000000011011111000011111011000;
        6'd08:obs<=32'b0000000111011101000010111011100;
        6'd09:obs<=32'b0000000111111101000010111011100;
        6'd10:obs<=32'b0000000101111101000010111111100;
        6'd11:obs<=32'b0000000111111111000011111111100;
        6'd12:obs<=32'b0000000111111111000011111111100;
        6'd13:obs<=32'b0000000111111111000011111111100;
        6'd14:obs<=32'b0000000011111111000011111111100;
        6'd15:obs<=32'b0000000011111111111111111111000;
        6'd16:obs<=32'b0000000001111000000000011111000;
        6'd17:obs<=32'b0000000001110000000000000111000;
        6'd18:obs<=32'b0000000001100000000000000111000;
        6'd19:obs<=32'b0000000010110000000000000101000;
        6'd20:obs<=32'b0000000011111000000000001111100;
        6'd21:obs<=32'b0000000011111111111111111111000;
        6'd22:obs<=32'b0000000001110111000011111111000;
        6'd23:obs<=32'b0000000001111111000011111011000;
        6'd24:obs<=32'b0000000001111111000011111011000;
        6'd25:obs<=32'b0000000001111111000011111011000;
        6'd26:obs<=32'b0000000001111111000011111011000;
        6'd27:obs<=32'b0000000001111111000011111111000;
        6'd28:obs<=32'b0000000011111111000011111111000;
        6'd29:obs<=32'b0000000011111111000011111011000;
        6'd30:obs<=32'b0000000001111111000011111011000;
        6'd31:obs<=32'b0000000001111111000011111011000;
        6'd32:obs<=32'b0000000001111111000011111111000;
        6'd33:obs<=32'b0000000011111111000011111111000;
        6'd34:obs<=32'b0000000101111111111111111111100;
        6'd35:obs<=32'b0000000101111000000110011111100;
        6'd36:obs<=32'b0000000101111000001110001111100;
        6'd37:obs<=32'b0000000111110000000000001111100;
        6'd38:obs<=32'b0000000111110000000000001111100;
        6'd39:obs<=32'b0000000111110000000000001111100;
        6'd40:obs<=32'b0000000111111111111111111111100;
        6'd41:obs<=32'b0000000011111111001011111111000;
        6'd42:obs<=32'b0000000001111111111111111111000;
        6'd43:obs<=32'b0000000001111111111111111111000;
        6'd44:obs<=32'b0000000001111111111111111110000;
        6'd45:obs<=32'b0000000001111111111111111110000;
        6'd46:obs<=32'b0000000000111111111111111100000;
        6'd47:obs<=32'b0000000000111111111111111100000;
        6'd48:obs<=32'b0000000000111111111111111100000;
        6'd49:obs<=32'b0000000000111111111111111100000;
    endcase
end
endmodule

module SCORE_DATA_DC(clk_25MHz,count,data,data_adrs,score_t);
input clk_25MHz;
input [4:0] data_adrs;
input [3:0] count;
output reg [0:19] data;
output reg [0:99] score_t;
always @(posedge clk_25MHz)
begin
    case(count)
    4'd0:
        begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000011000000000;
        5'd03:data<=20'b00000011111111000000;
        5'd04:data<=20'b00000111111111100000;
        5'd05:data<=20'b00001111111111110000;
        5'd06:data<=20'b00001111111111110000;
        5'd07:data<=20'b00011111000011111000;
        5'd08:data<=20'b00011110000011111000;
        5'd09:data<=20'b00011110000001111000;
        5'd10:data<=20'b00111110000001111000;
        5'd11:data<=20'b00111110000001111000;
        5'd12:data<=20'b00111110000001111100;
        5'd13:data<=20'b00111100000001111100;
        5'd14:data<=20'b00111100000001111100;
        5'd15:data<=20'b00111100000001111100;
        5'd16:data<=20'b00111100000001111100;
        5'd17:data<=20'b00111100000001111100;
        5'd18:data<=20'b00111100000001111100;
        5'd19:data<=20'b00111110000001111100;
        5'd20:data<=20'b00111110000001111000;
        5'd21:data<=20'b00111110000001111000;
        5'd22:data<=20'b00111110000001111000;
        5'd23:data<=20'b00111110000011111000;
        5'd24:data<=20'b00011111000011111000;
        5'd25:data<=20'b00011111100111110000;
        5'd26:data<=20'b00011111111111110000;
        5'd27:data<=20'b00001111111111100000;
        5'd28:data<=20'b00000111111111000000;
        5'd29:data<=20'b00000011111110000000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;    
        endcase
        end
    4'd1:begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000000000000000;
        5'd04:data<=20'b00000001111000000000;
        5'd05:data<=20'b00000011111000000000;
        5'd06:data<=20'b00000111111000000000;
        5'd07:data<=20'b00011111111000000000;
        5'd08:data<=20'b00011111111000000000;
        5'd09:data<=20'b00011101111000000000;
        5'd10:data<=20'b00011001111000000000;
        5'd11:data<=20'b00000001111000000000;
        5'd12:data<=20'b00000001111000000000;
        5'd13:data<=20'b00000001111000000000;
        5'd14:data<=20'b00000001111000000000;
        5'd15:data<=20'b00000001111000000000;
        5'd16:data<=20'b00000001111000000000;
        5'd17:data<=20'b00000001111000000000;
        5'd18:data<=20'b00000001111000000000;
        5'd19:data<=20'b00000001111000000000;
        5'd20:data<=20'b00000001111000000000;
        5'd21:data<=20'b00000001111000000000;
        5'd22:data<=20'b00000001111000000000;
        5'd23:data<=20'b00000001111000000000;
        5'd24:data<=20'b00000001111000000000;
        5'd25:data<=20'b00000001111100000000;
        5'd26:data<=20'b00011111111111100000;
        5'd27:data<=20'b00011111111111100000;
        5'd28:data<=20'b00011111111111100000;
        5'd29:data<=20'b00011111111111100000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
        end
    4'd2:
        begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000001111100000000;
        5'd03:data<=20'b00000111111111000000;
        5'd04:data<=20'b00011111111111100000;
        5'd05:data<=20'b00011111111111100000;
        5'd06:data<=20'b00011111111111110000;
        5'd07:data<=20'b00011100011111110000;
        5'd08:data<=20'b00011000001111110000;
        5'd09:data<=20'b00000000000111110000;
        5'd10:data<=20'b00000000000111110000;
        5'd11:data<=20'b00000000000111110000;
        5'd12:data<=20'b00000000000111110000;
        5'd13:data<=20'b00000000001111110000;
        5'd14:data<=20'b00000000001111100000;
        5'd15:data<=20'b00000000001111100000;
        5'd16:data<=20'b00000000011111000000;
        5'd17:data<=20'b00000000111111000000;
        5'd18:data<=20'b00000000111110000000;
        5'd19:data<=20'b00000001111100000000;
        5'd20:data<=20'b00000011111000000000;
        5'd21:data<=20'b00000111111000000000;
        5'd22:data<=20'b00001111110000000000;
        5'd23:data<=20'b00001111100000000000;
        5'd24:data<=20'b00011111000000000000;
        5'd25:data<=20'b00011111111111111000;
        5'd26:data<=20'b00111111111111111000;
        5'd27:data<=20'b00111111111111111000;
        5'd28:data<=20'b00011111111111111000;
        5'd29:data<=20'b00011111111111110000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
        end
    4'd3:
        begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000011000000000;
            5'd03:data<=20'b00000111111111000000;
            5'd04:data<=20'b00001111111111100000;
            5'd05:data<=20'b00011111111111100000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011100001111110000;
            5'd08:data<=20'b00010000000111110000;
            5'd09:data<=20'b00000000000111110000;
            5'd10:data<=20'b00000000000111110000;
            5'd11:data<=20'b00000000000111110000;
            5'd12:data<=20'b00000000000111110000;
            5'd13:data<=20'b00000000001111100000;
            5'd14:data<=20'b00000111111111000000;
            5'd15:data<=20'b00001111111110000000;
            5'd16:data<=20'b00001111111111000000;
            5'd17:data<=20'b00000111111111110000;
            5'd18:data<=20'b00000000011111110000;
            5'd19:data<=20'b00000000000111111000;
            5'd20:data<=20'b00000000000011111000;
            5'd21:data<=20'b00000000000011111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011111000;
            5'd24:data<=20'b00010000000111111000;
            5'd25:data<=20'b00111100001111111000;
            5'd26:data<=20'b00111111111111110000;
            5'd27:data<=20'b00111111111111100000;
            5'd28:data<=20'b00011111111111000000;
            5'd29:data<=20'b00001111111110000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
            endcase
        end
    4'd4:
    begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000011111100000;
        5'd04:data<=20'b00000000011111100000;
        5'd05:data<=20'b00000000111111100000;
        5'd06:data<=20'b00000000111111100000;
        5'd07:data<=20'b00000001111111100000;
        5'd08:data<=20'b00000001111111100000;
        5'd09:data<=20'b00000011110111100000;
        5'd10:data<=20'b00000011110111100000;
        5'd11:data<=20'b00000111100111100000;
        5'd12:data<=20'b00000111100111100000;
        5'd13:data<=20'b00001111000111100000;
        5'd14:data<=20'b00001111000111100000;
        5'd15:data<=20'b00011110000111100000;
        5'd16:data<=20'b00011110000111100000;
        5'd17:data<=20'b00111100000111100000;
        5'd18:data<=20'b00111100000111100000;
        5'd19:data<=20'b00111000000111100000;
        5'd20:data<=20'b00111111111111111100;
        5'd21:data<=20'b00111111111111111100;
        5'd22:data<=20'b00111111111111111100;
        5'd23:data<=20'b00111111111111111100;
        5'd24:data<=20'b00000000000111110000;
        5'd25:data<=20'b00000000000111100000;
        5'd26:data<=20'b00000000000111100000;
        5'd27:data<=20'b00000000000111100000;
        5'd28:data<=20'b00000000000111100000;
        5'd29:data<=20'b00000000000111100000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd5:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00001111111111100000;
            5'd04:data<=20'b00011111111111110000;
            5'd05:data<=20'b00011111111111110000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011111111111100000;
            5'd08:data<=20'b00011110000000000000;
            5'd09:data<=20'b00011110000000000000;
            5'd10:data<=20'b00011110000000000000;
            5'd11:data<=20'b00011110000000000000;
            5'd12:data<=20'b00011110000000000000;
            5'd13:data<=20'b00011111111100000000;
            5'd14:data<=20'b00011111111111000000;
            5'd15:data<=20'b00011111111111100000;
            5'd16:data<=20'b00011111111111110000;
            5'd17:data<=20'b00001100011111111000;
            5'd18:data<=20'b00000000000111111000;
            5'd19:data<=20'b00000000000011111000;
            5'd20:data<=20'b00000000000011111000;
            5'd21:data<=20'b00000000000011111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011111000;
            5'd24:data<=20'b00000000000111111000;
            5'd25:data<=20'b00011000001111110000;
            5'd26:data<=20'b00011111111111110000;
            5'd27:data<=20'b00011111111111100000;
            5'd28:data<=20'b00011111111111000000;
            5'd29:data<=20'b00001111111100000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd6:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00000000111111110000;
            5'd04:data<=20'b00000011111111110000;
            5'd05:data<=20'b00000011111111110000;
            5'd06:data<=20'b00000111111111110000;
            5'd07:data<=20'b00001111100000000000;
            5'd08:data<=20'b00001111000000000000;
            5'd09:data<=20'b00011111000000000000;
            5'd10:data<=20'b00011110000000000000;
            5'd11:data<=20'b00011110000000000000;
            5'd12:data<=20'b00011110000000000000;
            5'd13:data<=20'b00011110011111000000;
            5'd14:data<=20'b00011111111111110000;
            5'd15:data<=20'b00011111111111111000;
            5'd16:data<=20'b00111111111111111000;
            5'd17:data<=20'b00111111000011111100;
            5'd18:data<=20'b00111110000001111100;
            5'd19:data<=20'b00011110000001111100;
            5'd20:data<=20'b00011110000001111100;
            5'd21:data<=20'b00011110000001111100;
            5'd22:data<=20'b00011110000001111100;
            5'd23:data<=20'b00011110000001111100;
            5'd24:data<=20'b00011111000001111000;
            5'd25:data<=20'b00011111100011111000;
            5'd26:data<=20'b00001111111111111000;
            5'd27:data<=20'b00001111111111110000;
            5'd28:data<=20'b00000111111111100000;
            5'd29:data<=20'b00000001111110000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd7:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00011111111111111000;
            5'd04:data<=20'b00111111111111111000;
            5'd05:data<=20'b00111111111111111000;
            5'd06:data<=20'b00111111111111111000;
            5'd07:data<=20'b00011111111111111000;
            5'd08:data<=20'b00000000000011111000;
            5'd09:data<=20'b00000000000011111000;
            5'd10:data<=20'b00000000000111110000;
            5'd11:data<=20'b00000000000111110000;
            5'd12:data<=20'b00000000000111110000;
            5'd13:data<=20'b00000000001111100000;
            5'd14:data<=20'b00000000001111100000;
            5'd15:data<=20'b00000000001111000000;
            5'd16:data<=20'b00000000011111000000;
            5'd17:data<=20'b00000000011111000000;
            5'd18:data<=20'b00000000111110000000;
            5'd19:data<=20'b00000000111110000000;
            5'd20:data<=20'b00000000111110000000;
            5'd21:data<=20'b00000001111100000000;
            5'd22:data<=20'b00000001111100000000;
            5'd23:data<=20'b00000011111100000000;
            5'd24:data<=20'b00000011111000000000;
            5'd25:data<=20'b00000011111000000000;
            5'd26:data<=20'b00000111110000000000;
            5'd27:data<=20'b00000111110000000000;
            5'd28:data<=20'b00000111110000000000;
            5'd29:data<=20'b00000111100000000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd8:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000001000000000;
            5'd03:data<=20'b00000011111111000000;
            5'd04:data<=20'b00000111111111100000;
            5'd05:data<=20'b00001111111111110000;
            5'd06:data<=20'b00011111101111111000;
            5'd07:data<=20'b00011111000011111000;
            5'd08:data<=20'b00011110000001111000;
            5'd09:data<=20'b00011110000001111000;
            5'd10:data<=20'b00011110000001111000;
            5'd11:data<=20'b00011111000011111000;
            5'd12:data<=20'b00011111000111110000;
            5'd13:data<=20'b00001111111111100000;
            5'd14:data<=20'b00001111111111100000;
            5'd15:data<=20'b00000111111111000000;
            5'd16:data<=20'b00000011111111000000;
            5'd17:data<=20'b00000111111111110000;
            5'd18:data<=20'b00001111101111110000;
            5'd19:data<=20'b00011111000111111000;
            5'd20:data<=20'b00011110000011111000;
            5'd21:data<=20'b00111110000001111100;
            5'd22:data<=20'b00111100000001111100;
            5'd23:data<=20'b00111100000001111100;
            5'd24:data<=20'b00111110000001111000;
            5'd25:data<=20'b00111111000011111000;
            5'd26:data<=20'b00011111111111111000;
            5'd27:data<=20'b00011111111111110000;
            5'd28:data<=20'b00001111111111100000;
            5'd29:data<=20'b00000011111111000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd9:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000011000000000;
            5'd03:data<=20'b00000011111111000000;
            5'd04:data<=20'b00000111111111100000;
            5'd05:data<=20'b00001111111111110000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011111000011111000;
            5'd08:data<=20'b00111110000011111000;
            5'd09:data<=20'b00111110000001111000;
            5'd10:data<=20'b00111100000001111000;
            5'd11:data<=20'b00111100000001111000;
            5'd12:data<=20'b00111110000001111000;
            5'd13:data<=20'b00111110000001111000;
            5'd14:data<=20'b00111110000001111000;
            5'd15:data<=20'b00011111000111111000;
            5'd16:data<=20'b00011111111111111000;
            5'd17:data<=20'b00011111111111111000;
            5'd18:data<=20'b00001111111111111000;
            5'd19:data<=20'b00000011111001111000;
            5'd20:data<=20'b00000000000001111000;
            5'd21:data<=20'b00000000000001111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011110000;
            5'd24:data<=20'b00000000000111110000;
            5'd25:data<=20'b00011000001111100000;
            5'd26:data<=20'b00011111111111100000;
            5'd27:data<=20'b00011111111111000000;
            5'd28:data<=20'b00011111111110000000;
            5'd29:data<=20'b00001111111000000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd10:
    begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000000000000000;
        5'd04:data<=20'b00000000000000000000;
        5'd05:data<=20'b00000000000000000000;
        5'd06:data<=20'b00000000000000000000;
        5'd07:data<=20'b00000000000000000000;
        5'd08:data<=20'b00000000000000000000;
        5'd09:data<=20'b00000000000000000000;
        5'd10:data<=20'b00000000011111000000;
        5'd11:data<=20'b00000000011111000000;
        5'd12:data<=20'b00000000011111000000;
        5'd13:data<=20'b00000000011111000000;
        5'd14:data<=20'b00000000000000000000;
        5'd15:data<=20'b00000000000000000000;
        5'd16:data<=20'b00000000000000000000;
        5'd17:data<=20'b00000000000000000000;
        5'd18:data<=20'b00000000000000000000;
        5'd19:data<=20'b00000000000000000000;
        5'd20:data<=20'b00000000000000000000;
        5'd21:data<=20'b00000000000000000000;
        5'd22:data<=20'b00000000000000000000;
        5'd23:data<=20'b00000000011111000000;
        5'd24:data<=20'b00000000011111000000;
        5'd25:data<=20'b00000000011111000000;
        5'd26:data<=20'b00000000011111000000;
        5'd27:data<=20'b00000000000000000000;
        5'd28:data<=20'b00000000000000000000;
        5'd29:data<=20'b00000000000000000000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
    end
    default:
        data<=0;    
    endcase
end
always @(posedge clk_25MHz)
begin
    case(data_adrs)
        5'd00:score_t<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd01:score_t<=100'b0000000110000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000;
        5'd02:score_t<=100'b0000111111110000000000011111110000000000011111111100000000001111111110000000001111111111110000000000;
        5'd03:score_t<=100'b0001111111111000000001111111111100000000111111111110000000001111111111100000001111111111110000000000;
        5'd04:score_t<=100'b0011111111111000000011111111111110000001111111111111000000001111111111110000001111111111110000000000;
        5'd05:score_t<=100'b0011100000011000000011110000011110000011110000001111100000001110000011110000001111000000000000000000;
        5'd06:score_t<=100'b0111100000000000000111100000000110000111100000000011100000001110000001111000001110000000000000000000;
        5'd07:score_t<=100'b0111000000000000000111000000000000000111000000000011110000001110000001111000001110000000000000000000;
        5'd08:score_t<=100'b0111000000000000001111000000000000000111000000000001110000001110000000111000001110000000000000000000;
        5'd09:score_t<=100'b0111000000000000001110000000000000001111000000000001110000001110000000111000001110000000000000000000;
        5'd10:score_t<=100'b0111100000000000001110000000000000001110000000000001111000001110000000111000001110000000000000001100;
        5'd11:score_t<=100'b0111100000000000011110000000000000001110000000000000111000001110000000111000001110000000000000001110;
        5'd12:score_t<=100'b0011110000000000011100000000000000001110000000000000111000001110000001111000001110000000000000001110;
        5'd13:score_t<=100'b0011111000000000011100000000000000001110000000000000111000001110000001110000001110000000000000001110;
        5'd14:score_t<=100'b0001111110000000011100000000000000001110000000000000111000001110000111100000001111111111100000001110;
        5'd15:score_t<=100'b0000111111000000011100000000000000001110000000000000111000001111111111100000001111111111100000000000;
        5'd16:score_t<=100'b0000011111110000011100000000000000011110000000000000111000001111111110000000001111111111100000000000;
        5'd17:score_t<=100'b0000000111111000011100000000000000001110000000000000111000001111111111000000001111000000000000000000;
        5'd18:score_t<=100'b0000000011111000011100000000000000001110000000000000111000001110000111000000001110000000000000000000;
        5'd19:score_t<=100'b0000000000111100011100000000000000001110000000000000111000001110000011100000001110000000000000000000;
        5'd20:score_t<=100'b0000000000111100011100000000000000001110000000000000111000001110000011100000001110000000000000000000;
        5'd21:score_t<=100'b0000000000011100011110000000000000001110000000000001111000001110000001110000001110000000000000000000;
        5'd22:score_t<=100'b0000000000011100001110000000000000001110000000000001110000001110000001110000001110000000000000000000;
        5'd23:score_t<=100'b0000000000011100001110000000000000001111000000000001110000001110000001110000001110000000000000000000;
        5'd24:score_t<=100'b0000000000011100001111000000000000000111000000000011110000001110000001111000001110000000000000000000;
        5'd25:score_t<=100'b0000000000011100000111000000000010000111100000000011100000001110000000111000001110000000000000000000;
        5'd26:score_t<=100'b0110000000111000000111100000001110000111100000000111100000001110000000111000001110000000000000001110;
        5'd27:score_t<=100'b0111100001111000000011111000111110000011111000011111000000001110000000111100001111000000000000001110;
        5'd28:score_t<=100'b0111111111110000000011111111111100000001111111111110000000001110000000011100001111111111111000001110;
        5'd29:score_t<=100'b0011111111100000000001111111111000000000111111111100000000001110000000011100001111111111111000001110;
        5'd30:score_t<=100'b0001111111000000000000011111100000000000001111111000000000001110000000011100000111111111111000001110;
        5'd31:score_t<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
end
endmodule
