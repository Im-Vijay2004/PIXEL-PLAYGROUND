module PING_PONG(clk,clk_out,push11,push12,push21,push22,start,r,g,b,hcount,vcount,rst_pp);
    input clk,clk_out,rst_pp;
    output [3:0] r, g, b;
    input [9:0] hcount, vcount;
    wire clk_out2;//100mhz clock 
    wire [2:0]count_1,count_2;
    wire [4:0] score_adrs;
    wire [7:0] win_adrs;
    wire [0:149] score1,score2;
    wire [0:361] win;
    wire [1:0]playerwin;
    wire [9:0] paddle1_x , paddle1_y, paddle1_y2 ,paddle2_x ,paddle2_y,paddle2_y2 ,ball_x , ball_y ;     
    input push11, push12, push21, push22,start;
    
    
    SCORE_DATA_PP scoreone(clk_out,count_1,score1,score_adrs);
    SCORE_DATA_PP scoretwo(clk_out,count_2,score2,score_adrs);
    player_win_PP win1(clk_out,playerwin,win,win_adrs);
    clk_100hz_PP clk2(clk, clk_out2);
    disp_write_PP disp(clk_out,hcount,vcount,paddle1_x,paddle2_x,paddle1_y,paddle1_y2,paddle2_y,paddle2_y2,ball_x,ball_y,r,g,b,count1,score_adrs,score1,score2,win,win_adrs);
    paddle_movement_PP paddle(clk_out2,push11,push12,push21,push22,paddle1_y,paddle1_y2,paddle2_y,paddle2_y2,paddle1_x,paddle2_x);
    box_move_PP box(clk_out2,start,paddle1_y,paddle1_y2,paddle2_y,paddle2_y2,paddle1_x,paddle2_x,ball_x,ball_y,count_1,count_2,playerwin,rst_pp);

endmodule

`timescale 1ns / 1ps
module SCORE_DATA_PP(clk_25MHz,count, data, data_adrs);
    input clk_25MHz;
    input [4:0] data_adrs;
    input [2:0] count;
    output reg [0:149] data;

    always @(posedge clk_25MHz) begin
        case(count)
            3'd0: begin
                case(data_adrs)
        5'd00:data<=150'b00000000000111111100000000000111111100000000000000000000000000011111110000000000011111110000000000000000000000000000111111100000000000111111100000000000;
        5'd01:data<=150'b00000000011111111111000000011111111111000000000000000000000001111111111100000001111111111100000000000000000000000011111111111000000011111111111000000000;
        5'd02:data<=150'b00000000111111111111100000111111111111100000000000000000000011111111111111000011111111111110000000000000000000000111111111111100000111111111111100000000;
        5'd03:data<=150'b00000001111111111111110011111111111111110000000000000000000111111111111111100111111111111111000000000000000000001111111111111110011111111111111110000000;
        5'd04:data<=150'b00000011111111111111111111111111111111110000000000000000000111111111111111111111111111111111100000000000000000011111111111111111111111111111111110000000;
        5'd05:data<=150'b00000011111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000000000000011111111111111111111111111111111111000000;
        5'd06:data<=150'b00000111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111000000;
        5'd07:data<=150'b00000111111111111111111111111111111111111100000000000000011111111111111111111111111111111111110000000000000000111111111111111111111111111111111111100000;
        5'd08:data<=150'b00000111111111111111111111111111111111111100000000000000011111111111111111111111111111111111110000000000000000111111111111111111111111111111111111100000;
        5'd09:data<=150'b00000111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111000000000000000111111111111111111111111111111111111100000;
        5'd10:data<=150'b00000111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111000000000000000111111111111111111111111111111111111100000;
        5'd11:data<=150'b00000111111111111111111111111111111111111100000000000000011111111111111111111111111111111111110000000000000000111111111111111111111111111111111111100000;
        5'd12:data<=150'b00000111111111111111111111111111111111111100000000000000011111111111111111111111111111111111110000000000000000111111111111111111111111111111111111100000;
        5'd13:data<=150'b00000111111111111111111111111111111111111100000000000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111000000;
        5'd14:data<=150'b00000011111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000000000000011111111111111111111111111111111111000000;
        5'd15:data<=150'b00000011111111111111111111111111111111111000000000000000001111111111111111111111111111111111100000000000000000011111111111111111111111111111111111000000;
        5'd16:data<=150'b00000011111111111111111111111111111111110000000000000000000111111111111111111111111111111111100000000000000000011111111111111111111111111111111110000000;
        5'd17:data<=150'b00000001111111111111111111111111111111100000000000000000000011111111111111111111111111111111000000000000000000001111111111111111111111111111111100000000;
        5'd18:data<=150'b00000000111111111111111111111111111111100000000000000000000001111111111111111111111111111110000000000000000000000111111111111111111111111111111100000000;
        5'd19:data<=150'b00000000011111111111111111111111111111000000000000000000000001111111111111111111111111111100000000000000000000000011111111111111111111111111111000000000;
        5'd20:data<=150'b00000000001111111111111111111111111110000000000000000000000000111111111111111111111111111100000000000000000000000011111111111111111111111111110000000000;
        5'd21:data<=150'b00000000001111111111111111111111111100000000000000000000000000011111111111111111111111111000000000000000000000000001111111111111111111111111100000000000;
        5'd22:data<=150'b00000000000111111111111111111111111000000000000000000000000000001111111111111111111111110000000000000000000000000000111111111111111111111111000000000000;
        5'd23:data<=150'b00000000000011111111111111111111111000000000000000000000000000000111111111111111111111100000000000000000000000000000011111111111111111111110000000000000;
        5'd24:data<=150'b00000000000001111111111111111111110000000000000000000000000000000011111111111111111111000000000000000000000000000000001111111111111111111100000000000000;
        5'd25:data<=150'b00000000000000111111111111111111000000000000000000000000000000000001111111111111111110000000000000000000000000000000000111111111111111111000000000000000;
        5'd26:data<=150'b00000000000000011111111111111110000000000000000000000000000000000000111111111111111100000000000000000000000000000000000011111111111111110000000000000000;
        5'd27:data<=150'b00000000000000000111111111111100000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000111111111111100000000000000000;
        5'd28:data<=150'b00000000000000000011111111111000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000011111111111000000000000000000;
        5'd29:data<=150'b00000000000000000001111111100000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000001111111100000000000000000000;
        5'd30:data<=150'b00000000000000000000011111000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000011111000000000000000000000;
        5'd31:data<=150'b00000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000;
      
                    default: data <= 150'b0;
                endcase
            end
            3'd1: begin
                case(data_adrs)
        5'd00:data<=150'b0000000000011111110000000000011111110000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000;
        5'd01:data<=150'b0000000001111111111100000001111111111100000000000000000000000111111111110000000111111111110000000000000000000000000000000000000000000000000000000000000;
        5'd02:data<=150'b0000000011111111111110000011111111111110000000000000000000001111111111111100001111111111111000000000000000000000000000000000000000000000000000000000000;
        5'd03:data<=150'b0000000111111111111111001111111111111111000000000000000000011111111111111110011111111111111100000000000000000000000000000000000000000000000000000000000;
        5'd04:data<=150'b0000001111111111111111111111111111111111000000000000000000011111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
        5'd05:data<=150'b0000001111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
        5'd06:data<=150'b0000011111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
        5'd07:data<=150'b0000011111111111111111111111111111111111110000000000000001111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
        5'd08:data<=150'b0000011111111111111111111111111111111111110000000000000001111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
        5'd09:data<=150'b0000011111111111111111111111111111111111110000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000;
        5'd10:data<=150'b0000011111111111111111111111111111111111110000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000;
        5'd11:data<=150'b0000011111111111111111111111111111111111110000000000000001111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
        5'd12:data<=150'b0000011111111111111111111111111111111111110000000000000001111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
        5'd13:data<=150'b0000011111111111111111111111111111111111110000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
        5'd14:data<=150'b0000001111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
        5'd15:data<=150'b0000001111111111111111111111111111111111100000000000000000111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
        5'd16:data<=150'b0000001111111111111111111111111111111111000000000000000000011111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
        5'd17:data<=150'b0000000111111111111111111111111111111110000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
        5'd18:data<=150'b0000000011111111111111111111111111111110000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
        5'd19:data<=150'b0000000001111111111111111111111111111100000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
        5'd20:data<=150'b0000000000111111111111111111111111111000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
        5'd21:data<=150'b0000000000111111111111111111111111110000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000;
        5'd22:data<=150'b0000000000011111111111111111111111100000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
        5'd23:data<=150'b0000000000001111111111111111111111100000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000;
        5'd24:data<=150'b0000000000000111111111111111111111000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000;
        5'd25:data<=150'b0000000000000011111111111111111100000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000;
        5'd26:data<=150'b0000000000000001111111111111111000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000;
        5'd27:data<=150'b0000000000000000011111111111110000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000;
        5'd28:data<=150'b0000000000000000001111111111100000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000;
        5'd29:data<=150'b0000000000000000000111111110000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000;
        5'd30:data<=150'b0000000000000000000001111100000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd31:data<=150'b0000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000;
                  
            default: data <= 150'b0;
        endcase
        end
        3'd2: begin
                case(data_adrs)
        5'd00:data<=150'b0000000000011111110000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd01:data<=150'b0000000001111111111100000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd02:data<=150'b0000000011111111111110000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd03:data<=150'b0000000111111111111111001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd04:data<=150'b0000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd05:data<=150'b0000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd06:data<=150'b0000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd07:data<=150'b0000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd08:data<=150'b0000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd09:data<=150'b0000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd10:data<=150'b0000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd11:data<=150'b0000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd12:data<=150'b0000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd13:data<=150'b0000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd14:data<=150'b0000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd15:data<=150'b0000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd16:data<=150'b0000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd17:data<=150'b0000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd18:data<=150'b0000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd19:data<=150'b0000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd20:data<=150'b0000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd21:data<=150'b0000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd22:data<=150'b0000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd23:data<=150'b0000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd24:data<=150'b0000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd25:data<=150'b0000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd26:data<=150'b0000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd27:data<=150'b0000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd28:data<=150'b0000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd29:data<=150'b0000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd30:data<=150'b0000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd31:data<=150'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        default: data <= 150'b0; 
        endcase        
            
            end
        default: data <= 0;
        endcase
    end
endmodule


module player_win_PP(clk_25MHz,player,win,data_adrs);
input clk_25MHz;
input [7:0] data_adrs;
input [1:0]player;
output reg [0:361]win;


always @(posedge clk_25MHz) begin
   case(player)
    3'd1: begin
          case(data_adrs)
8'd000:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd001:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd002:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd003:win<=362'b0000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd004:win<=362'b0011111111111111111111111111111110000000000000000000000011111111111110000000000000000000000000000000000000000000000000111111111111110000000000000001111111111111100000000000000000000000011111111111111000000011111111111111111111111111111111111111110000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000;
8'd005:win<=362'b0011111111111111111111111111111111110000000000000000000011111111111110000000000000000000000000000000000000000000000001111111111111110000000000000000111111111111110000000000000000000000011111111111111000000011111111111111111111111111111111111111110000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000001111111111100;
8'd006:win<=362'b0011111111111111111111111111111111111100000000000000000011111111111110000000000000000000000000000000000000000000000001111111111111110000000000000000111111111111110000000000000000000000111111111111110000000011111111111111111111111111111111111111110000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000011111111111110;
8'd007:win<=362'b0011111111111111111111111111111111111111000000000000000011111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111000000000000000000000111111111111110000000011111111111111111111111111111111111111110000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000111111111111110;
8'd008:win<=362'b0011111111111111111111111111111111111111100000000000000011111111111110000000000000000000000000000000000000000000000011111111111111111000000000000000011111111111111000000000000000000001111111111111100000000011111111111111111111111111111111111111110000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111110;
8'd009:win<=362'b0011111111111111111111111111111111111111110000000000000011111111111110000000000000000000000000000000000000000000000011111111111111111000000000000000001111111111111100000000000000000001111111111111100000000011111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111000000000000000000000000000000000000000000000011111111111111110;
8'd010:win<=362'b0011111111111111111111111111111111111111111000000000000011111111111110000000000000000000000000000000000000000000000011111111111111111100000000000000001111111111111100000000000000000011111111111111000000000011111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111100000000000000000000000000000000000000000000111111111111111110;
8'd011:win<=362'b0011111111111111111111111111111111111111111100000000000011111111111110000000000000000000000000000000000000000000000111111111111111111100000000000000000111111111111110000000000000000011111111111110000000000011111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111110000000000000000000000000000000000000000011111111111111111110;
8'd012:win<=362'b0011111111111111111111111111111111111111111110000000000011111111111110000000000000000000000000000000000000000000000111111111111111111110000000000000000111111111111110000000000000000111111111111110000000000011111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111110000000000000000000000000000000000000001111111111111111111110;
8'd013:win<=362'b0011111111111111111111111111111111111111111110000000000011111111111110000000000000000000000000000000000000000000001111111111111111111110000000000000000011111111111111000000000000000111111111111100000000000011111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111111111110;
8'd014:win<=362'b0011111111111110000000000000111111111111111111000000000011111111111110000000000000000000000000000000000000000000001111111111111111111110000000000000000011111111111111000000000000001111111111111100000000000011111111111110000000000000000000000000000000000000011111111111110000000000001111111111111111111000000000000000000000000000000000111111111111111111111111110;
8'd015:win<=362'b0011111111111110000000000000001111111111111111000000000011111111111110000000000000000000000000000000000000000000001111111111111111111111000000000000000001111111111111100000000000001111111111111000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000001111111111111111000000000000000000000000000000011111111111111111111111111110;
8'd016:win<=362'b0011111111111110000000000000000011111111111111000000000011111111111110000000000000000000000000000000000000000000011111111111111111111111000000000000000001111111111111100000000000011111111111111000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000011111111111111000000000000000000000000000000011111111111111111111111111110;
8'd017:win<=362'b0011111111111110000000000000000011111111111111100000000011111111111110000000000000000000000000000000000000000000011111111111111111111111000000000000000000111111111111110000000000011111111111110000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000011111111111111100000000000000000000000000000011111111111111111111111111110;
8'd018:win<=362'b0011111111111110000000000000000001111111111111100000000011111111111110000000000000000000000000000000000000000000011111111111011111111111100000000000000000011111111111110000000000111111111111110000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000001111111111111100000000000000000000000000000011111111111111111111111111110;
8'd019:win<=362'b0011111111111110000000000000000001111111111111100000000011111111111110000000000000000000000000000000000000000000111111111111011111111111100000000000000000011111111111111000000000111111111111100000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000001111111111111100000000000000000000000000000011111111111111111111111111110;
8'd020:win<=362'b0011111111111110000000000000000000111111111111100000000011111111111110000000000000000000000000000000000000000000111111111111001111111111100000000000000000001111111111111000000001111111111111100000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000001111111111111100000000000000000000000000000011111111111111011111111111110;
8'd021:win<=362'b0011111111111110000000000000000000111111111111100000000011111111111110000000000000000000000000000000000000000000111111111110001111111111110000000000000000001111111111111100000001111111111111000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000001111111111111100000000000000000000000000000011111111111110011111111111110;
8'd022:win<=362'b0011111111111110000000000000000000111111111111100000000011111111111110000000000000000000000000000000000000000001111111111110001111111111110000000000000000000111111111111100000011111111111111000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000001111111111111000000000000000000000000000000011111111111000011111111111110;
8'd023:win<=362'b0011111111111110000000000000000000111111111111100000000011111111111110000000000000000000000000000000000000000001111111111110000111111111111000000000000000000111111111111110000011111111111110000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000001111111111111000000000000000000000000000000011111111110000011111111111110;
8'd024:win<=362'b0011111111111110000000000000000000111111111111100000000011111111111110000000000000000000000000000000000000000011111111111100000111111111111000000000000000000011111111111110000111111111111100000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000001111111111111000000000000000000000000000000011111111000000011111111111110;
8'd025:win<=362'b0011111111111110000000000000000000111111111111100000000011111111111110000000000000000000000000000000000000000011111111111100000111111111111000000000000000000011111111111111000111111111111100000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000001111111111111000000000000000000000000000000011111000000000011111111111110;
8'd026:win<=362'b0011111111111110000000000000000001111111111111100000000011111111111110000000000000000000000000000000000000000011111111111100000011111111111100000000000000000001111111111111001111111111111000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000011111111111110000000000000000000000000000000000000000000000011111111111110;
8'd027:win<=362'b0011111111111110000000000000000001111111111111100000000011111111111110000000000000000000000000000000000000000111111111111000000011111111111100000000000000000001111111111111101111111111111000000000000000000011111111111111111111111111111111111110000000000000011111111111110000000000000000111111111111110000000000000000000000000000000000000000000000011111111111110;
8'd028:win<=362'b0011111111111110000000000000000011111111111111000000000011111111111110000000000000000000000000000000000000000111111111111000000011111111111100000000000000000000111111111111111111111111110000000000000000000011111111111111111111111111111111111110000000000000011111111111110000000000000001111111111111100000000000000000000000000000000000000000000000011111111111110;
8'd029:win<=362'b0011111111111110000000000000000111111111111111000000000011111111111110000000000000000000000000000000000000000111111111111000000001111111111110000000000000000000011111111111111111111111110000000000000000000011111111111111111111111111111111111110000000000000011111111111110000000000011111111111111111100000000000000000000000000000000000000000000000011111111111110;
8'd030:win<=362'b0011111111111110000000000000011111111111111111000000000011111111111110000000000000000000000000000000000000001111111111110000000001111111111110000000000000000000011111111111111111111111100000000000000000000011111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011111111111110;
8'd031:win<=362'b0011111111111111011111111111111111111111111110000000000011111111111110000000000000000000000000000000000000001111111111110000000001111111111110000000000000000000001111111111111111111111100000000000000000000011111111111111111111111111111111111110000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111110;
8'd032:win<=362'b0011111111111111111111111111111111111111111110000000000011111111111110000000000000000000000000000000000000001111111111110000000000111111111111000000000000000000001111111111111111111111000000000000000000000011111111111111111111111111111111111110000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011111111111110;
8'd033:win<=362'b0011111111111111111111111111111111111111111100000000000011111111111110000000000000000000000000000000000000011111111111100000000000111111111111000000000000000000000111111111111111111111000000000000000000000011111111111111111111111111111111111110000000000000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000011111111111110;
8'd034:win<=362'b0011111111111111111111111111111111111111111000000000000011111111111110000000000000000000000000000000000000011111111111100000000000111111111111000000000000000000000111111111111111111110000000000000000000000011111111111111111111111111111111111110000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111110;
8'd035:win<=362'b0011111111111111111111111111111111111111111000000000000011111111111110000000000000000000000000000000000000011111111111100000000000011111111111100000000000000000000011111111111111111110000000000000000000000011111111111111111111111111111111111110000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111110;
8'd036:win<=362'b0011111111111111111111111111111111111111110000000000000011111111111110000000000000000000000000000000000000111111111111000000000000011111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111111111111111111111111000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000011111111111110;
8'd037:win<=362'b0011111111111111111111111111111111111111100000000000000011111111111110000000000000000000000000000000000000111111111111000000000000011111111111110000000000000000000001111111111111111000000000000000000000000011111111111111111111111111111111111110000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011111111111110;
8'd038:win<=362'b0011111111111111111111111111111111111110000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000001111111111110000000000000000000001111111111111111000000000000000000000000011111111111110000000000000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111110;
8'd039:win<=362'b0011111111111111111111111111111111111000000000000000000011111111111110000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000111111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011111111111110;
8'd040:win<=362'b0011111111111111111111111111111111100000000000000000000011111111111110000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000111111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111111000000000011111111111111111000000000000000000000000000000000000000000000000011111111111110;
8'd041:win<=362'b0011111111111111111111111111111000000000000000000000000011111111111110000000000000000000000000000000000011111111111111111111111111111111111111111000000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000011111111111111100000000000000000000000000000000000000000000000011111111111110;
8'd042:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111110000000000000000000000000000000000011111111111111111111111111111111111111111000000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000111111111111110000000000000000000000000000000000000000000000011111111111110;
8'd043:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111110000000000000000000000000000000000011111111111111111111111111111111111111111100000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000111111111111110000000000000000000000000000000000000000000000011111111111110;
8'd044:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111110000000000000000000000000000000000111111111111111111111111111111111111111111100000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000011111111111110000000000000000000000000000000000000000000000011111111111110;
8'd045:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111110000000000000000000000000000000000111111111111111111111111111111111111111111100000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000001111111111111000000000000000000000000000000000000000000000011111111111110;
8'd046:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111110000000000000000000000000000000000111111111111111111111111111111111111111111110000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000001111111111111000000000000000000000000000000000000000000000011111111111110;
8'd047:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111110000000000000000000000000000000001111111111111111111111111111111111111111111110000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000001111111111111000000000000000000000000000000000000000000000011111111111110;
8'd048:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111110000000000000000000000000000000001111111111111111111111111111111111111111111111000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000000111111111111100000000000000000000000000000000000000000000011111111111110;
8'd049:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111110000000000000000000000000000000001111111111111111111111111111111111111111111111000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000000111111111111100000000000000000000000000000000000000000000011111111111110;
8'd050:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111110000000000000000000000000000000011111111111110000000000000000000001111111111111000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000000111111111111100000000000000000000000000000000000000000000011111111111110;
8'd051:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111111111111111111111111111110000000011111111111110000000000000000000000111111111111100000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000000111111111111100000000000000000000000000000000000000000000011111111111110;
8'd052:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111000000111111111111110000000000000000000000111111111111100000000000000000011111111111110000000000000000000000000011111111111111111111111111111111111111110000000000011111111111110000000000000000000011111111111110000000000000000000000000000000000000000000011111111111110;
8'd053:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111000000111111111111100000000000000000000000111111111111100000000000000000011111111111110000000000000000000000000011111111111111111111111111111111111111110000000000011111111111110000000000000000000011111111111110000000000000000000000000000000000000000000011111111111110;
8'd054:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111000000111111111111100000000000000000000000011111111111110000000000000000011111111111110000000000000000000000000011111111111111111111111111111111111111110000000000011111111111110000000000000000000011111111111110000000000000000000000000000000000000000000011111111111110;
8'd055:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111000001111111111111100000000000000000000000011111111111110000000000000000011111111111110000000000000000000000000011111111111111111111111111111111111111110000000000011111111111110000000000000000000011111111111111000000000000000000000000000000000000000000011111111111110;
8'd056:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111000001111111111111000000000000000000000000011111111111110000000000000000011111111111110000000000000000000000000011111111111111111111111111111111111111110000000000011111111111110000000000000000000001111111111111000000000000000000000000000000000000000000011111111111110;
8'd057:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111000001111111111111000000000000000000000000001111111111111000000000000000011111111111110000000000000000000000000011111111111111111111111111111111111111110000000000011111111111110000000000000000000001111111111111000000000000000000000000000000000000000000011111111111110;
8'd058:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111000011111111111111000000000000000000000000001111111111111000000000000000011111111111110000000000000000000000000011111111111111111111111111111111111111110000000000011111111111110000000000000000000001111111111111000000000000000000000000000000000000000000011111111111110;
8'd059:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111000011111111111110000000000000000000000000001111111111111000000000000000011111111111110000000000000000000000000011111111111111111111111111111111111111110000000000011111111111110000000000000000000001111111111111100000000000000000000000000000000000000000011111111111110;
8'd060:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111000011111111111110000000000000000000000000001111111111111100000000000000011111111111110000000000000000000000000011111111111111111111111111111111111111110000000000011111111111110000000000000000000000111111111111100000000000000000000000000000000000000000011111111111110;
8'd061:win<=362'b0011111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111000111111111111110000000000000000000000000000111111111111100000000000000011111111111110000000000000000000000000011111111111111111111111111111111111111110000000000011111111111110000000000000000000000111111111111100000000000000000000000000000000000000000011111111111110;
8'd062:win<=362'b0001111111111110000000000000000000000000000000000000000001111111111111111111111111111111111111000111111111111100000000000000000000000000000111111111111100000000000000011111111111110000000000000000000000000011111111111111111111111111111111111111110000000000011111111111110000000000000000000000111111111111100000000000000000000000000000000000000000011111111111100;
8'd063:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd064:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd065:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd066:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd067:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd068:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd069:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd070:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd071:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd072:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd073:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd074:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd075:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd076:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd077:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd078:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd079:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd080:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd081:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd082:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd083:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd084:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd085:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd086:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd087:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd088:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd089:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd090:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd091:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd092:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd093:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd094:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd095:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd096:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd097:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd098:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd099:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd100:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd101:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd102:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd103:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd104:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000001111111111111100000000000000000000001111111111111000000011111111111100000000000000111111111111100000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd105:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000001111111111111100000000000000000000011111111111111000000011111111111110000000000000111111111111110000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd106:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000001111111111111100000000000000000000011111111111110000000011111111111110000000000000111111111111110000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd107:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000001111111111111100000000000000000000011111111111110000000011111111111110000000000000111111111111111000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd108:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000011111111111111110000000000000000000011111111111110000000011111111111110000000000000111111111111111100000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd109:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000011111111111111110000000000000000000111111111111100000000011111111111110000000000000111111111111111100000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd110:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000011111111111111110000000000000000000111111111111100000000011111111111110000000000000111111111111111110000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd111:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000111111111111111110000000000000000000111111111111100000000011111111111110000000000000111111111111111111000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd112:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000111111111111111111000000000000000000111111111111000000000011111111111110000000000000111111111111111111000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd113:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000111111111111111111000000000000000001111111111111000000000011111111111110000000000000111111111111111111100000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd114:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000111111111111111111000000000000000001111111111111000000000011111111111110000000000000111111111111111111110000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd115:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000001111111111111111111100000000000000001111111111111000000000011111111111110000000000000111111111111111111110000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd116:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000001111111111111111111100000000000000001111111111110000000000011111111111110000000000000111111111111111111111000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd117:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000001111111111111111111100000000000000011111111111110000000000011111111111110000000000000111111111111111111111100000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd118:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000001111111111111111111100000000000000011111111111110000000000011111111111110000000000000111111111111111111111100000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd119:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000011111111111111111111110000000000000011111111111100000000000011111111111110000000000000111111111111111111111110000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd120:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000011111111111111111111110000000000000011111111111100000000000011111111111110000000000000111111111111111111111111000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd121:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000011111111111111111111110000000000000111111111111100000000000011111111111110000000000000111111111111111111111111000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd122:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000011111111110111111111110000000000000111111111111000000000000011111111111110000000000000111111111111111111111111100000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd123:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000111111111110011111111111000000000000111111111111000000000000011111111111110000000000000111111111111111111111111110000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd124:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000111111111110011111111111000000000000111111111111000000000000011111111111110000000000000111111111111111111111111111000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd125:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000111111111110011111111111000000000001111111111111000000000000011111111111110000000000000111111111111011111111111111000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd126:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000001111111111100011111111111000000000001111111111110000000000000011111111111110000000000000111111111111001111111111111100000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd127:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000001111111111100001111111111100000000001111111111110000000000000011111111111110000000000000111111111111001111111111111110000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd128:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000001111111111100001111111111100000000001111111111110000000000000011111111111110000000000000111111111111000111111111111110000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd129:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000001111111111000001111111111100000000011111111111100000000000000011111111111110000000000000111111111111000011111111111111000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd130:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000011111111111000001111111111110000000011111111111100000000000000011111111111110000000000000111111111111000011111111111111100000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd131:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000011111111111000000111111111110000000011111111111100000000000000011111111111110000000000000111111111111000001111111111111100000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd132:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000011111111111000000111111111110000000111111111111000000000000000011111111111110000000000000111111111111000000111111111111110000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd133:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000011111111110000000111111111110000000111111111111000000000000000011111111111110000000000000111111111111000000111111111111111000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd134:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111110000000011111111111000000111111111111000000000000000011111111111110000000000000111111111111000000011111111111111000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd135:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111110000000011111111111000000111111111111000000000000000011111111111110000000000000111111111111000000001111111111111100000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd136:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000111111111110000000011111111111000001111111111110000000000000000011111111111110000000000000111111111111000000001111111111111110000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd137:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000111111111100000000011111111111000001111111111110000000000000000011111111111110000000000000111111111111000000000111111111111110000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd138:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100001111111111100000000001111111111100001111111111110000000000000000011111111111110000000000000111111111111000000000011111111111111000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd139:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100001111111111100000000001111111111100001111111111100000000000000000011111111111110000000000000111111111111000000000011111111111111100111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd140:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110001111111111100000000001111111111100011111111111100000000000000000011111111111110000000000000111111111111000000000001111111111111100111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd141:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110011111111111000000000001111111111110011111111111100000000000000000011111111111110000000000000111111111111000000000000111111111111110111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd142:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110011111111111000000000000111111111110011111111111000000000000000000011111111111110000000000000111111111111000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd143:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110011111111111000000000000111111111110011111111111000000000000000000011111111111110000000000000111111111111000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd144:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111011111111111000000000000111111111110111111111111000000000000000000011111111111110000000000000111111111111000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd145:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000111111111111111111111111000000000000000000011111111111110000000000000111111111111000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd146:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000011111111111111111111110000000000000000000011111111111110000000000000111111111111000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd147:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000011111111111111111111110000000000000000000011111111111110000000000000111111111111000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd148:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000011111111111111111111110000000000000000000011111111111110000000000000111111111111000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd149:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000011111111111111111111100000000000000000000011111111111110000000000000111111111111000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd150:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000001111111111111111111100000000000000000000011111111111110000000000000111111111111000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd151:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000001111111111111111111100000000000000000000011111111111110000000000000111111111111000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd152:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000001111111111111111111100000000000000000000011111111111110000000000000111111111111000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd153:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000111111111111111111000000000000000000000011111111111110000000000000111111111111000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd154:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000111111111111111111000000000000000000000011111111111110000000000000111111111111000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd155:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000111111111111111111000000000000000000000011111111111110000000000000111111111111000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd156:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111111111111111110000000000000000000000011111111111110000000000000111111111111000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd157:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000011111111111111110000000000000000000000011111111111110000000000000111111111111000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd158:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000011111111111111110000000000000000000000011111111111110000000000000111111111111000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd159:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000011111111111111100000000000000000000000011111111111110000000000000111111111111000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd160:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000011111111111111100000000000000000000000011111111111110000000000000111111111111000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd161:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000001111111111111100000000000000000000000011111111111110000000000000111111111111000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd162:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000001111111111111000000000000000000000000011111111111100000000000000111111111111000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd163:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd164:win<=362'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
default:win <= 362'b0;
endcase
end 

    3'd2: begin
        case(data_adrs)
8'd000:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd001:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd002:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd003:win<=362'b00111111111111111111111111111110000000000000000000000011111111111100000000000000000000000000000000000000000000000111111111111100000000000000011111111111111000000000000000000000001111111111111100000011111111111111111111111111111111111111100000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd004:win<=362'b00111111111111111111111111111111110000000000000000000011111111111100000000000000000000000000000000000000000000000111111111111110000000000000011111111111111000000000000000000000011111111111111000000011111111111111111111111111111111111111100000000001111111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111110000000000000000000;
8'd005:win<=362'b00111111111111111111111111111111111100000000000000000011111111111100000000000000000000000000000000000000000000001111111111111110000000000000001111111111111100000000000000000000011111111111111000000011111111111111111111111111111111111111100000000001111111111111111111111111111111111110000000000000000000000000000000000000000000011111111111111111110000000000000000;
8'd006:win<=362'b00111111111111111111111111111111111111000000000000000011111111111100000000000000000000000000000000000000000000001111111111111110000000000000000111111111111100000000000000000000111111111111110000000011111111111111111111111111111111111111100000000001111111111111111111111111111111111111100000000000000000000000000000000000000001111111111111111111111000000000000000;
8'd007:win<=362'b00111111111111111111111111111111111111100000000000000011111111111100000000000000000000000000000000000000000000001111111111111111000000000000000111111111111110000000000000000000111111111111110000000011111111111111111111111111111111111111100000000001111111111111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000;
8'd008:win<=362'b00111111111111111111111111111111111111110000000000000011111111111100000000000000000000000000000000000000000000011111111111111111000000000000000011111111111110000000000000000001111111111111100000000011111111111111111111111111111111111111100000000001111111111111111111111111111111111111111000000000000000000000000000000000001111111111111111111111111111000000000000;
8'd009:win<=362'b00111111111111111111111111111111111111111000000000000011111111111100000000000000000000000000000000000000000000011111111111111111000000000000000011111111111111000000000000000001111111111111100000000011111111111111111111111111111111111111100000000001111111111111111111111111111111111111111100000000000000000000000000000000011111111111111111111111111111100000000000;
8'd010:win<=362'b00111111111111111111111111111111111111111100000000000011111111111100000000000000000000000000000000000000000000111111111111111111100000000000000001111111111111000000000000000011111111111111000000000011111111111111111111111111111111111111100000000001111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000;
8'd011:win<=362'b00111111111111111111111111111111111111111100000000000011111111111100000000000000000000000000000000000000000000111111111111111111100000000000000001111111111111100000000000000011111111111111000000000011111111111111111111111111111111111111100000000001111111111111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111110000000000;
8'd012:win<=362'b00111111111111111111111111111111111111111110000000000011111111111100000000000000000000000000000000000000000000111111111111111111110000000000000000111111111111100000000000000111111111111110000000000011111111111111111111111111111111111111100000000001111111111111111111111111111111111111111110000000000000000000000000000001111111111111111111111111111111111000000000;
8'd013:win<=362'b00111111111111000000000000111111111111111110000000000011111111111100000000000000000000000000000000000000000001111111111111111111110000000000000000111111111111110000000000000111111111111100000000000011111111111110000000000000000000000000000000000001111111111111000000000001111111111111111111000000000000000000000000000001111111111111111111111111111111111000000000;
8'd014:win<=362'b00111111111111000000000000000111111111111111000000000011111111111100000000000000000000000000000000000000000001111111111111111111110000000000000000011111111111110000000000000111111111111100000000000011111111111110000000000000000000000000000000000001111111111111000000000000001111111111111111000000000000000000000000000011111111111111100000011111111111111100000000;
8'd015:win<=362'b00111111111111000000000000000011111111111111000000000011111111111100000000000000000000000000000000000000000001111111111111111111111000000000000000011111111111111000000000001111111111111000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000011111111111111000000000000000000000000000011111111111110000000001111111111111100000000;
8'd016:win<=362'b00111111111111000000000000000001111111111111000000000011111111111100000000000000000000000000000000000000000011111111111111111111111000000000000000001111111111111000000000001111111111111000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000001111111111111000000000000000000000000000011111111111100000000000111111111111100000000;
8'd017:win<=362'b00111111111111000000000000000001111111111111100000000011111111111100000000000000000000000000000000000000000011111111111011111111111000000000000000001111111111111100000000011111111111110000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000001111111111111000000000000000000000000000011111111111100000000000011111111111110000000;
8'd018:win<=362'b00111111111111000000000000000000111111111111100000000011111111111100000000000000000000000000000000000000000011111111111011111111111100000000000000000111111111111100000000011111111111110000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000001111111111111000000000000000000000000000111111111111000000000000011111111111110000000;
8'd019:win<=362'b00111111111111000000000000000000111111111111100000000011111111111100000000000000000000000000000000000000000111111111111001111111111100000000000000000011111111111110000000111111111111100000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000001111111111111000000000000000000000000000111111111111000000000000011111111111110000000;
8'd020:win<=362'b00111111111111000000000000000000111111111111100000000011111111111100000000000000000000000000000000000000000111111111110001111111111100000000000000000011111111111110000000111111111111100000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000000111111111111000000000000000000000000000111111111111000000000000001111111111110000000;
8'd021:win<=362'b00111111111111000000000000000000111111111111100000000011111111111100000000000000000000000000000000000000001111111111110001111111111110000000000000000001111111111111000001111111111111000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000001111111111111000000000000000000000000000111111111110000000000000001111111111110000000;
8'd022:win<=362'b00111111111111000000000000000000111111111111100000000011111111111100000000000000000000000000000000000000001111111111110000111111111110000000000000000001111111111111000001111111111111000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000001111111111111000000000000000000000000000111111111110000000000000001111111111110000000;
8'd023:win<=362'b00111111111111000000000000000000111111111111100000000011111111111100000000000000000000000000000000000000001111111111100000111111111111000000000000000000111111111111100011111111111110000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000001111111111111000000000000000000000000000011111111110000000000000011111111111110000000;
8'd024:win<=362'b00111111111111000000000000000000111111111111100000000011111111111100000000000000000000000000000000000000011111111111100000111111111111000000000000000000111111111111100011111111111100000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000001111111111110000000000000000000000000000000000000000000000000000011111111111100000000;
8'd025:win<=362'b00111111111111000000000000000001111111111111100000000011111111111100000000000000000000000000000000000000011111111111100000011111111111000000000000000000011111111111110111111111111100000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000011111111111110000000000000000000000000000000000000000000000000000011111111111100000000;
8'd026:win<=362'b00111111111111000000000000000001111111111111000000000011111111111100000000000000000000000000000000000000011111111111000000011111111111100000000000000000011111111111111111111111111000000000000000000011111111111111111111111111111111111100000000000001111111111111000000000000000111111111111100000000000000000000000000000000000000000000000000000111111111111100000000;
8'd027:win<=362'b00111111111111000000000000000011111111111111000000000011111111111100000000000000000000000000000000000000111111111111000000011111111111100000000000000000001111111111111111111111111000000000000000000011111111111111111111111111111111111100000000000001111111111111000000000000011111111111111100000000000000000000000000000000000000000000000000000111111111111100000000;
8'd028:win<=362'b00111111111111000000000000000111111111111111000000000011111111111100000000000000000000000000000000000000111111111111000000001111111111100000000000000000001111111111111111111111110000000000000000000011111111111111111111111111111111111100000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000001111111111111000000000;
8'd029:win<=362'b00111111111111100000000000111111111111111110000000000011111111111100000000000000000000000000000000000000111111111110000000001111111111110000000000000000000111111111111111111111110000000000000000000011111111111111111111111111111111111100000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111000000000;
8'd030:win<=362'b00111111111111111111111111111111111111111110000000000011111111111100000000000000000000000000000000000001111111111110000000001111111111110000000000000000000111111111111111111111100000000000000000000011111111111111111111111111111111111100000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111110000000000;
8'd031:win<=362'b00111111111111111111111111111111111111111100000000000011111111111100000000000000000000000000000000000001111111111110000000000111111111110000000000000000000011111111111111111111100000000000000000000011111111111111111111111111111111111100000000000001111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111110000000000;
8'd032:win<=362'b00111111111111111111111111111111111111111100000000000011111111111100000000000000000000000000000000000001111111111100000000000111111111111000000000000000000001111111111111111111000000000000000000000011111111111111111111111111111111111100000000000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000001111111111111100000000000;
8'd033:win<=362'b00111111111111111111111111111111111111111000000000000011111111111100000000000000000000000000000000000011111111111100000000000111111111111000000000000000000001111111111111111111000000000000000000000011111111111111111111111111111111111100000000000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111111000000000000;
8'd034:win<=362'b00111111111111111111111111111111111111110000000000000011111111111100000000000000000000000000000000000011111111111100000000000011111111111000000000000000000000111111111111111110000000000000000000000011111111111111111111111111111111111100000000000001111111111111111111111111111111111110000000000000000000000000000000000000000000000000000111111111111110000000000000;
8'd035:win<=362'b00111111111111111111111111111111111111100000000000000011111111111100000000000000000000000000000000000111111111111000000000000011111111111100000000000000000000111111111111111110000000000000000000000011111111111111111111111111111111111100000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000001111111111111100000000000000;
8'd036:win<=362'b00111111111111111111111111111111111111000000000000000011111111111100000000000000000000000000000000000111111111111000000000000011111111111100000000000000000000011111111111111100000000000000000000000011111111111110000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000011111111111111000000000000000;
8'd037:win<=362'b00111111111111111111111111111111111100000000000000000011111111111100000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000011111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111111111110000000000000000;
8'd038:win<=362'b00111111111111111111111111111111100000000000000000000011111111111100000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000011111111111111100000000000000000;
8'd039:win<=362'b00111111111111111111111111111100000000000000000000000011111111111100000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000011111111111111100000000000000000000000000000000000000000111111111111111000000000000000000;
8'd040:win<=362'b00111111111111000000000000000000000000000000000000000011111111111100000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000111111111111100000000000000000000000000000000000000001111111111111110000000000000000000;
8'd041:win<=362'b00111111111111000000000000000000000000000000000000000011111111111100000000000000000000000000000000011111111111111111111111111111111111111111000000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000011111111111110000000000000000000000000000000000000011111111111111100000000000000000000;
8'd042:win<=362'b00111111111111000000000000000000000000000000000000000011111111111100000000000000000000000000000000011111111111111111111111111111111111111111000000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000011111111111110000000000000000000000000000000000000111111111111111000000000000000000000;
8'd043:win<=362'b00111111111111000000000000000000000000000000000000000011111111111100000000000000000000000000000000011111111111111111111111111111111111111111100000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000001111111111110000000000000000000000000000000000001111111111111110000000000000000000000;
8'd044:win<=362'b00111111111111000000000000000000000000000000000000000011111111111100000000000000000000000000000000111111111111111111111111111111111111111111100000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000001111111111111000000000000000000000000000000000011111111111111100000000000000000000000;
8'd045:win<=362'b00111111111111000000000000000000000000000000000000000011111111111100000000000000000000000000000000111111111111111111111111111111111111111111100000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000001111111111111000000000000000000000000000000000111111111111111000000000000000000000000;
8'd046:win<=362'b00111111111111000000000000000000000000000000000000000011111111111100000000000000000000000000000000111111111111111111111111111111111111111111110000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000000111111111111000000000000000000000000000000001111111111111110000000000000000000000000;
8'd047:win<=362'b00111111111111000000000000000000000000000000000000000011111111111100000000000000000000000000000001111111111111111111111111111111111111111111110000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000000111111111111100000000000000000000000000000011111111111111000000000000000000000000000;
8'd048:win<=362'b00111111111111000000000000000000000000000000000000000011111111111110000000000000000000000000000001111111111111000000000000000000001111111111111000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000000111111111111100000000000000000000000000001111111111111110000000000000000000000000000;
8'd049:win<=362'b00111111111111000000000000000000000000000000000000000011111111111111111111111111111111111100000011111111111110000000000000000000001111111111111000000000000000001111111111111000000000000000000000000011111111111110000000000000000000000000000000000001111111111111000000000000000000111111111111100000000000000000000000000011111111111111100000000000000000000000000000;
8'd050:win<=362'b00111111111111000000000000000000000000000000000000000011111111111111111111111111111111111100000011111111111110000000000000000000000111111111111000000000000000001111111111111000000000000000000000000011111111111111111111111111111111111111100000000001111111111111000000000000000000011111111111100000000000000000000000000111111111111111111111111111111111111111000000;
8'd051:win<=362'b00111111111111000000000000000000000000000000000000000011111111111111111111111111111111111100000011111111111100000000000000000000000111111111111100000000000000001111111111111000000000000000000000000011111111111111111111111111111111111111100000000001111111111111000000000000000000011111111111110000000000000000000000001111111111111111111111111111111111111111000000;
8'd052:win<=362'b00111111111111000000000000000000000000000000000000000011111111111111111111111111111111111100000111111111111100000000000000000000000111111111111100000000000000001111111111111000000000000000000000000011111111111111111111111111111111111111100000000001111111111111000000000000000000011111111111110000000000000000000000001111111111111111111111111111111111111111000000;
8'd053:win<=362'b00111111111111000000000000000000000000000000000000000011111111111111111111111111111111111100000111111111111100000000000000000000000111111111111100000000000000001111111111111000000000000000000000000011111111111111111111111111111111111111100000000001111111111111000000000000000000011111111111110000000000000000000000001111111111111111111111111111111111111111000000;
8'd054:win<=362'b00111111111111000000000000000000000000000000000000000011111111111111111111111111111111111100000111111111111100000000000000000000000011111111111110000000000000001111111111111000000000000000000000000011111111111111111111111111111111111111100000000001111111111111000000000000000000001111111111111000000000000000000000001111111111111111111111111111111111111111000000;
8'd055:win<=362'b00111111111111000000000000000000000000000000000000000011111111111111111111111111111111111100001111111111111000000000000000000000000011111111111110000000000000001111111111111000000000000000000000000011111111111111111111111111111111111111100000000001111111111111000000000000000000001111111111111000000000000000000000001111111111111111111111111111111111111111000000;
8'd056:win<=362'b00111111111111000000000000000000000000000000000000000011111111111111111111111111111111111100001111111111111000000000000000000000000011111111111110000000000000001111111111111000000000000000000000000011111111111111111111111111111111111111100000000001111111111111000000000000000000001111111111111000000000000000000000001111111111111111111111111111111111111111000000;
8'd057:win<=362'b00111111111111000000000000000000000000000000000000000011111111111111111111111111111111111100001111111111111000000000000000000000000001111111111111000000000000001111111111111000000000000000000000000011111111111111111111111111111111111111100000000001111111111111000000000000000000001111111111111000000000000000000000001111111111111111111111111111111111111111000000;
8'd058:win<=362'b00111111111111000000000000000000000000000000000000000011111111111111111111111111111111111100011111111111110000000000000000000000000001111111111111000000000000001111111111111000000000000000000000000011111111111111111111111111111111111111100000000001111111111111000000000000000000000111111111111100000000000000000000011111111111111111111111111111111111111111000000;
8'd059:win<=362'b00111111111111000000000000000000000000000000000000000011111111111111111111111111111111111100011111111111110000000000000000000000000001111111111111000000000000001111111111111000000000000000000000000011111111111111111111111111111111111111100000000001111111111111000000000000000000000111111111111100000000000000000000001111111111111111111111111111111111111111000000;
8'd060:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd061:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd062:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd063:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd064:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd065:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd066:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd067:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd068:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd069:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd070:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd071:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd072:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd073:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd074:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd075:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd076:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd077:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd078:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd079:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd080:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd081:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd082:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd083:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd084:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd085:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd086:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd087:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd088:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd089:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd090:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd091:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd092:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000111111111110000000000000000000000011111111111000000001111111111100000000000000111111111110000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd093:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000001111111111111000000000000000000000111111111111100000011111111111110000000000000111111111111000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd094:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000001111111111111000000000000000000000111111111111000000011111111111110000000000000111111111111100000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd095:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000011111111111111100000000000000000001111111111111000000011111111111110000000000000111111111111110000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd096:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000011111111111111100000000000000000001111111111111000000011111111111110000000000000111111111111110000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd097:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000011111111111111100000000000000000001111111111111000000011111111111110000000000000111111111111111000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd098:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000011111111111111100000000000000000001111111111110000000011111111111110000000000000111111111111111100000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd099:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000111111111111111110000000000000000011111111111110000000011111111111110000000000000111111111111111110000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd100:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000111111111111111110000000000000000011111111111110000000011111111111110000000000000111111111111111110000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd101:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000111111111111111110000000000000000011111111111100000000011111111111110000000000000111111111111111111000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd102:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000111111111111111110000000000000000011111111111100000000011111111111110000000000000111111111111111111100000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd103:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000001111111111111111111000000000000000111111111111100000000011111111111110000000000000111111111111111111100000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd104:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000001111111111111111111000000000000000111111111111000000000011111111111110000000000000111111111111111111110000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd105:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000001111111111111111111000000000000000111111111111000000000011111111111110000000000000111111111111111111111000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd106:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000011111111111111111111000000000000000111111111111000000000011111111111110000000000000111111111111111111111000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd107:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000011111111111111111111100000000000001111111111111000000000011111111111110000000000000111111111111111111111100000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd108:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000011111111111111111111100000000000001111111111110000000000011111111111110000000000000111111111111111111111110000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd109:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000011111111111111111111100000000000001111111111110000000000011111111111110000000000000111111111111111111111110000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd110:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000111111111110111111111110000000000001111111111110000000000011111111111110000000000000111111111111111111111111000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd111:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000111111111110111111111110000000000011111111111100000000000011111111111110000000000000111111111111111111111111100000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd112:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000111111111100111111111110000000000011111111111100000000000011111111111110000000000000111111111111111111111111100000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd113:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000111111111100011111111110000000000011111111111100000000000011111111111110000000000000111111111110111111111111110000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd114:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000001111111111100011111111111000000000011111111111100000000000011111111111110000000000000111111111110011111111111111000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd115:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000001111111111100011111111111000000000111111111111000000000000011111111111110000000000000111111111110011111111111111000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd116:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000001111111111000011111111111000000000111111111111000000000000011111111111110000000000000111111111110001111111111111100000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd117:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000001111111111000001111111111000000000111111111111000000000000011111111111110000000000000111111111110000111111111111110000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd118:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000011111111111000001111111111100000000111111111110000000000000011111111111110000000000000111111111110000011111111111111000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd119:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000011111111111000001111111111100000001111111111110000000000000011111111111110000000000000111111111110000011111111111111000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd120:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000011111111110000001111111111100000001111111111110000000000000011111111111110000000000000111111111110000001111111111111100000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd121:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111110000000111111111110000001111111111100000000000000011111111111110000000000000111111111110000000111111111111110000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd122:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000111111111110000000111111111110000001111111111100000000000000011111111111110000000000000111111111110000000111111111111110000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd123:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000111111111100000000111111111110000011111111111100000000000000011111111111110000000000000111111111110000000011111111111111000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd124:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000111111111100000000111111111110000011111111111100000000000000011111111111110000000000000111111111110000000001111111111111100011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd125:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100001111111111100000000011111111111000011111111111000000000000000011111111111110000000000000111111111110000000001111111111111100011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd126:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100001111111111100000000011111111111000111111111111000000000000000011111111111110000000000000111111111110000000000111111111111110011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd127:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110001111111111000000000011111111111000111111111111000000000000000011111111111110000000000000111111111110000000000011111111111111011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd128:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110001111111111000000000011111111111000111111111110000000000000000011111111111110000000000000111111111110000000000011111111111111011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd129:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110011111111111000000000001111111111100111111111110000000000000000011111111111110000000000000111111111110000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd130:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110011111111111000000000001111111111101111111111110000000000000000011111111111110000000000000111111111110000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd131:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111011111111110000000000001111111111101111111111100000000000000000011111111111110000000000000111111111110000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd132:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000001111111111101111111111100000000000000000011111111111110000000000000111111111110000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd133:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000111111111111111111111100000000000000000011111111111110000000000000111111111110000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd134:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000111111111111111111111100000000000000000011111111111110000000000000111111111110000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd135:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000111111111111111111111000000000000000000011111111111110000000000000111111111110000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd136:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000011111111111111111111000000000000000000011111111111110000000000000111111111110000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd137:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000011111111111111111111000000000000000000011111111111110000000000000111111111110000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd138:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000011111111111111111110000000000000000000011111111111110000000000000111111111110000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd139:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000011111111111111111110000000000000000000011111111111110000000000000111111111110000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd140:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000001111111111111111110000000000000000000011111111111110000000000000111111111110000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd141:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000001111111111111111100000000000000000000011111111111110000000000000111111111110000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd142:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000001111111111111111100000000000000000000011111111111110000000000000111111111110000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd143:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000001111111111111111100000000000000000000011111111111110000000000000111111111110000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd144:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000111111111111111100000000000000000000011111111111110000000000000111111111110000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd145:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000111111111111111000000000000000000000011111111111110000000000000111111111110000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd146:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000111111111111111000000000000000000000011111111111110000000000000111111111110000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd147:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000111111111111111000000000000000000000011111111111110000000000000111111111110000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd148:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000011111111111110000000000000000000000011111111111110000000000000111111111110000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd149:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000011111111111110000000000000000000000001111111111110000000000000111111111110000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd150:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd151:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd152:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd153:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd154:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd155:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd156:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd157:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd158:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd159:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd160:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd161:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd162:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd163:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
8'd164:win<=362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
default: win <= 362'b0;
endcase 
end 
default: win <= 362'b0;
endcase
end 
endmodule


module clk_100hz_PP(clk_in,clk_out);
input clk_in;
output reg clk_out=0;
integer i;
always @(posedge clk_in)
begin
    if(i==499999)
    begin
        clk_out<=~clk_out;
        i<=0;
    end
    else
        i<=i+1;
end
endmodule

module disp_write_PP(clk,hcount,vcount,paddle1_x,paddle2_x,paddle1_y,paddle1_y2,paddle2_y,paddle2_y2,ball_x,ball_y,red,green,blue,count1,score_adrs,score1,score2,win,win_adrs);
input clk;
input [3:0]count1 = 4'b0001;
output reg [3:0] red, green, blue;
input [9:0] hcount, vcount;
input [9:0] paddle1_x,paddle2_x,paddle1_y,paddle1_y2,paddle2_y,paddle2_y2,ball_x,ball_y;
output reg [4:0] score_adrs;
output reg [7:0] win_adrs;
input [0:361] win;
input [0:149] score1,score2;
always @(posedge clk) begin
        if ((hcount >= 144 && hcount <= 784) && (vcount >= 35 && vcount <= 521)) 
        begin
            score_adrs <= vcount - 40;
            win_adrs <= vcount - 190;
           if ((hcount >= 620 && hcount <= 770) && (vcount > 40 && vcount < 72) && (score1[hcount - 620] == 1))
                {red, green, blue} <= {4'b0000, 4'b0000, 4'b1111};
           else if ((hcount >= 150 && hcount <= 300) && (vcount > 40 && vcount < 72) && (score2[hcount - 150] == 1))
                {red, green, blue} <= {4'b1111, 4'b0000, 4'b0000}; // Blue pixel for score
           else if ((hcount >= 280 && hcount <= 642) && (vcount > 190 && vcount < 355) && (win[hcount - 280] == 1))
                {red, green, blue} <= {4'b0110, 4'b0010, 4'b1111};
           else if ((hcount >= ball_x && hcount <= ball_x + 60) && (vcount >= ball_y && vcount <= ball_y + 60))
                {red, green, blue} <= {4'b0000, 4'b1111, 4'b0000}; // Ball: Green
            else if ((hcount >= paddle1_x && hcount <= paddle1_x + 30) && 
                     (vcount >= paddle1_y && vcount <= paddle1_y + 90))
                {red, green, blue} <= {4'b1111, 4'b0000, 4'b0000}; // Paddle 1: Red
            else if ((hcount >= paddle2_x && hcount <= paddle2_x + 30) && 
                     (vcount >= paddle2_y && vcount <= paddle2_y + 90))
                {red, green, blue} <= {4'b0000, 4'b0000, 4'b1111}; // Paddle 2: Blue
            else if ((hcount >= 454 && hcount <= 474))
                {red, green, blue} <= {4'b1111, 4'b1111, 4'b1111}; // Divider
            else
                {red, green, blue} <= {4'b0000, 4'b0000, 4'b0000}; // Background: White
        end else begin
            {red, green, blue} <= {4'b0000, 4'b0000, 4'b0000}; // Outside boundary: Black
        end
    end
endmodule

module paddle_movement_PP(clk_out2,push11,push12,push21,push22,paddle1_y,paddle1_y2,paddle2_y,paddle2_y2,paddle1_x,paddle2_x);
input clk_out2,push11,push12,push21,push22;
output reg [9:0]paddle1_x = 144,
             paddle1_y = 245,
             paddle1_y2 = 335,
             paddle2_x = 754,
             paddle2_y = 245,
             paddle2_y2 = 335;
             
 always @(posedge clk_out2) begin
        if (push11 && (paddle1_y2 < 521)) begin
            paddle1_y <= paddle1_y + 1;
            paddle1_y2 <= paddle1_y2 + 1;
        end else if (push12 && (paddle1_y > 35) ) begin
            paddle1_y <= paddle1_y - 1;
            paddle1_y2 <= paddle1_y2 - 1;
        end 
        else begin
             paddle1_y <= paddle1_y;
            paddle1_y2 <= paddle1_y2;
        end 
        
        
         if (push21 && (paddle2_y2 < 521) ) begin
            paddle2_y <= paddle2_y + 1;
            paddle2_y2 <= paddle2_y2 + 1;
        end else if (push22 && (paddle2_y > 35)) begin
            paddle2_y <= paddle2_y - 1;
            paddle2_y2 <= paddle2_y2 - 1;
        end 
        else begin
            paddle2_y <= paddle2_y;
            paddle2_y2 <= paddle2_y2;
        end
        
    end
endmodule

module box_move_PP(clk_out2, start, paddle1_y, paddle1_y2, paddle2_y, paddle2_y2, 
                paddle1_x, paddle2_x, ball_x, ball_y, count_1, count_2,playerwin,rst_pp);
    
    reg game_reset, game_start;
    input clk_out2, start,rst_pp;
    input [9:0] paddle1_y, paddle1_y2, paddle2_y, paddle2_y2, paddle1_x, paddle2_x;
    output reg [9:0] ball_x = 444, ball_y = 235;
    reg horizontal_dir, vertical_dir;
    reg [3:0] random_value = 4'b1011;
    reg [3:0] random_value1 = 4'b1011;
    output reg [2:0] count_1, count_2;
    output reg [1:0]playerwin;
    always @(posedge clk_out2) begin
        // Generate randomness continuously
        
        
        if (game_reset|rst_pp) begin
            // Reset game parameters
            
            ball_x <= 434;
            ball_y <= 245;
            game_start <= 0; 
            game_reset <= 0;
        end 
        else if (start && !game_start) begin
            game_start <= 1;
            count_1 <= 0;
            count_2 <= 0;
            playerwin <= 0; 
        end

        if (game_start) begin
            // Ball movement logic
            if ((ball_x + 50 >= paddle2_x && ball_x <= paddle2_x + 30) &&
                (ball_y + 50 >= paddle2_y && ball_y <= paddle2_y2)) begin
                horizontal_dir <= 0;
                random_value <= {random_value[2:0], random_value[3] ^ random_value[2]}; 
                vertical_dir <= random_value[0];
               
            end 
            else if ((ball_x <= paddle1_x + 30 && ball_x >= paddle1_x) &&
                     (ball_y + 50 >= paddle1_y && ball_y <= paddle1_y2)) begin
                horizontal_dir <= 1;
                random_value1 <= {random_value1[2:0], random_value1[3] ^ random_value1[2]}; 
                vertical_dir <= random_value1[0];
            end 
            
            // Randomize vertical movement periodically
            

            // Vertical boundary collision
            if (ball_y + 50 >= 521)
                vertical_dir <= 0;
            else if (ball_y <= 35)
                vertical_dir <= 1;

            // Update ball position
            if (horizontal_dir)
                ball_x <= ball_x + 1;
            else
                ball_x <= ball_x - 1;

            if (vertical_dir)
                ball_y <= ball_y + 1;
            else
                ball_y <= ball_y - 1;

            // Scoring logic
            if (ball_x <= 144) begin
                ball_x <= 464;
                ball_y <= 278;
                count_2 <= count_2 + 1;
            end 
            else if (ball_x + 50 >= 784) begin
                ball_x <= 464;
                ball_y <= 278;
                count_1 <= count_1 + 1;
            end

            // Game reset condition
            if ((count_1 <= 7 && count_1 > 2) || (count_2 <= 7 && count_2 > 2)) begin
                game_reset <= 1;
                if(count_1 > count_2)
                    playerwin <= 1;
                 else if(count_2> count_1) 
                    playerwin <= 2;
                 else 
                    playerwin <= 0;  
                
            end
        end
    end
endmodule
