`timescale 1ns / 1ps
module TIC_TAC_TOE(sys_clk,clk_25M,lt,rt,up,dn,reset1,enter,hcount,vcount,red,green,blue,win,rst_ttt);
input sys_clk,clk_25M,enter,reset1,rst_ttt;
input lt,rt,up,dn;
input [9:0] hcount,vcount;
output [1:0]win;
output [3:0] red,green,blue;
wire [9:0] select_x,select_y;
wire clk_1M;
wire [6:0]data_adrs;
wire [0:119]data;
wire [5:0] title_adrs;
wire [0:423] title;
wire [0:219] player;
wire [6:0] player_adrs;
wire [6:0] win_adrs;
wire [0:219] win1;
wire [1:0]sp0,sp1,sp2,sp3,sp4,sp5,sp6,sp7,sp8,data_sel;
//assign win=win_temp;
wire reset;
assign reset=reset1|rst_ttt;
CLK_10Hz Clk_div(sys_clk,clk_1M);
DATA_TTT bit(clk_25M,data,data_adrs,data_sel);
Title_TTT title_data(clk_25M,title,title_adrs,player,player_adrs);
WIN_LOGIC Winner(clk_25M,win1,win_adrs,win);
win game_end(clk_25M,sp0,sp1,sp2,sp3,sp4,sp5,sp6,sp7,sp8,win,reset);
DISP_WRITE_TTT Disp_w(clk_25M,hcount,vcount,red,green,blue,select_x,select_y,data_adrs,data,data_sel,title,title_adrs,player,player_adrs,win1,win_adrs,sp0,sp1,sp2,sp3,sp4,sp5,sp6,sp7,sp8);
game_fsm fsm(clk_1M,reset,up,dn,rt,lt,select_x,select_y,enter,sp0,sp1,sp2,sp3,sp4,sp5,sp6,sp7,sp8,win);
endmodule

module DISP_WRITE_TTT(clk_25M,hcount,vcount,red,green,blue,select_x,select_y,data_adrs,data,data_sel,title,title_adrs,player,player_adrs,win1,win_adrs,sp0,sp1,sp2,sp3,sp4,sp5,sp6,sp7,sp8);
input clk_25M;
input [9:0] hcount,vcount,select_x,select_y;
output reg [3:0] red,green,blue;
output reg [6:0] data_adrs;
input [0:119] data;
input [0:423] title;
input [0:219] player;
input [0:219] win1;
output reg [6:0] player_adrs;
output reg [5:0] title_adrs;
output reg [1:0]data_sel;
output reg [6:0] win_adrs;
input [1:0]sp0,sp1,sp2,sp3,sp4,sp5,sp6,sp7,sp8;
parameter   hmin=144,
            hmax=784,
            vmin=35,
            vmax=515;
parameter   box_h1=379,
            box_v1=108,
            box_h2=510,
            box_h3=640,
            box_v2=238,
            box_v3=368
;
always @(posedge clk_25M)
begin
    if((hcount>=hmin && hcount<=hmax) && (vcount>=vmin && vcount<=vmax))
        begin
            title_adrs<=vcount-40;
            player_adrs<=vcount-140;
            win_adrs<=vcount-250;
            if((hcount>=369 && hcount<=770) && (vcount>=98 && vcount<=500 ))
            begin
                
                 if((hcount>= box_h1 && hcount<=box_h1+119) && (vcount>=box_v1 && vcount<=box_v1+119 ))
                begin
                data_adrs=vcount-box_v1;
                data_sel=sp0;
                if(data[hcount-box_h1]==1)
                    {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                else if((hcount>= select_x && hcount<=select_x+119) && (vcount>=select_y && vcount<=select_y+119 ))
                begin
                    {red,green,blue}<={4'b0011,4'b1101,4'b1101};
                end
                else
                    {red,green,blue}<={4'b0011,4'b1101,4'b0100};
                end
                else if((hcount>= box_h2 && hcount<=box_h2+119) && (vcount>=box_v1 && vcount<=box_v1+119 ))
                begin
                data_adrs=vcount-box_v1;
                data_sel=sp1;
                if(data[hcount-box_h2]==1)
                    {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                else if((hcount>= select_x && hcount<=select_x+119) && (vcount>=select_y && vcount<=select_y+119 ))
                begin
                    {red,green,blue}<={4'b0011,4'b1101,4'b1101};
                end
                else
                    {red,green,blue}<={4'b0011,4'b1101,4'b0100};
                end
               
                else if((hcount>= box_h3 && hcount<=box_h3+119) && (vcount>=box_v1 && vcount<=box_v1+119 ))
                begin
                data_adrs=vcount-box_v1;
                data_sel=sp2;
                if(data[hcount-box_h3]==1)
                    {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                   else if((hcount>= select_x && hcount<=select_x+119) && (vcount>=select_y && vcount<=select_y+119 ))
                begin
                    {red,green,blue}<={4'b0011,4'b1101,4'b1101};
                end
                else
                    {red,green,blue}<={4'b0011,4'b1101,4'b0100};
                end
                
                else if((hcount>= box_h1 && hcount<=box_h1+119) && (vcount>=box_v2 && vcount<=box_v2+119 ))
                begin
                data_adrs=vcount-box_v2;
                data_sel=sp3;
                if(data[hcount-box_h1]==1)
                    {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                   else if((hcount>= select_x && hcount<=select_x+119) && (vcount>=select_y && vcount<=select_y+119 ))
                begin
                    {red,green,blue}<={4'b0011,4'b1101,4'b1101};
                end
                else
                    {red,green,blue}<={4'b0011,4'b1101,4'b0100};
                end
               
                else if((hcount>= box_h2 && hcount<=box_h2+119) && (vcount>=box_v2 && vcount<=box_v2+119 ))
                begin
                data_adrs=vcount-box_v2;
                data_sel=sp4;
                 if(data[hcount-box_h2-5]==1)
                    {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                  else if((hcount>= select_x && hcount<=select_x+119) && (vcount>=select_y && vcount<=select_y+119 ))
               begin
                    {red,green,blue}<={4'b0011,4'b1101,4'b1101};
                end
                else
                    {red,green,blue}<={4'b0011,4'b1101,4'b0100};
                end
                else if((hcount>= box_h3 && hcount<=box_h3+119) && (vcount>=box_v2 && vcount<=box_v2+119 ))
                begin
                data_adrs=vcount-box_v2;
                data_sel=sp5;
                if(data[hcount-box_h3+5]==1)
                    {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                else if((hcount>= select_x && hcount<=select_x+119) && (vcount>=select_y && vcount<=select_y+119 ))
                begin
                    {red,green,blue}<={4'b0011,4'b1101,4'b1101};
                end
                else
                    {red,green,blue}<={4'b0011,4'b1101,4'b0100};
                end
                else if((hcount>= box_h1 && hcount<=box_h1+119) && (vcount>=box_v3 && vcount<=box_v3+119 ))
                begin
                data_adrs=vcount-box_v3;
                data_sel=sp6;
                if(data[hcount-box_h1]==1)
                    {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                   else if((hcount>= select_x && hcount<=select_x+119) && (vcount>=select_y && vcount<=select_y+119 ))
                begin
                    {red,green,blue}<={4'b0011,4'b1101,4'b1101};
                end
                else
                    {red,green,blue}<={4'b0011,4'b1101,4'b0100};
                end
                else if((hcount>= box_h2 && hcount<=box_h2+119) && (vcount>=box_v3 && vcount<=box_v3+119 ))
                begin
                data_adrs=vcount-box_v3;
                data_sel=sp7;
                if(data[hcount-box_h2]==1)
                    {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                  else if((hcount>= select_x && hcount<=select_x+119) && (vcount>=select_y && vcount<=select_y+119 ))
                begin
                    {red,green,blue}<={4'b0011,4'b1101,4'b1101};
                end
                else
                    {red,green,blue}<={4'b0011,4'b1101,4'b0100};
                end
                else if((hcount>= box_h3 && hcount<=box_h3+119) && (vcount>=box_v3 && vcount<=box_v3+119 ))
                begin
                data_adrs=vcount-box_v3;
                data_sel=sp8;
                if(data[hcount-box_h1]==1)
                    {red,green,blue}<={4'b1111,4'b1111,4'b1111};
                       else if((hcount>= select_x && hcount<=select_x+119) && (vcount>=select_y && vcount<=select_y+119 ))
                begin
                    {red,green,blue}<={4'b0011,4'b1101,4'b1101};
                end
                else
                    {red,green,blue}<={4'b0011,4'b1101,4'b0100};
                end
                else
                    {red,green,blue}<={4'b0001,4'b0010,4'b0100}; //PLAY AREA BACKGROUND BROWN
            end
            else if((hcount>252 && hcount<676)&& (vcount>=40 && vcount<95)&& title[hcount-252]==1)
            begin
                {red,green,blue}<={4'b1111,4'b0101,4'b0111};
            end
            else if((hcount>=148 && hcount<367)&& (vcount>=140 && vcount<222)&& player[hcount-148]==1)
            begin
                {red,green,blue}<={4'b1111,4'b1111,4'b1111};
            end
            else if((hcount>=148 && hcount<367)&& (vcount>=250 && vcount<378)&& win1[hcount-148]==1)
            begin
                {red,green,blue}<={4'b0110,4'b0001,4'b0100};
            end
            else
            {red,green,blue}<={4'b0001,4'b0010,4'b0011};// ENTIRE BACKGROUND 
        end
    else
        begin
            {red,green,blue}<={4'b0000,4'b0000,4'b0000};   
        end
end
endmodule

module win(sys_clk,sp0,sp1,sp2,sp3,sp4,sp5,sp6,sp7,sp8,win,reset);
input [1:0]sp0,sp1,sp2,sp3,sp4,sp5,sp6,sp7,sp8;
input sys_clk,reset;
output reg [1:0]win;
always @(posedge sys_clk)
begin
if(reset)
begin 
    win<=0;
end 
else
begin
    if((sp0==1 && sp1==1 && sp2==1)||(sp3==1 && sp4==1 && sp5==1)||( sp6==1 && sp7==1 && sp8==1)||(sp0==1 && sp3==1 && sp6==1)||
    (sp1==1 && sp4==1 && sp7==1)||(sp2==1 && sp5==1 && sp8==1)||(sp0===1 && sp4==1 && sp8==1)||(sp2==1 && sp4==1 && sp6==1))
        win=2'b01;
    else if((sp0==2 && sp1==2 && sp2==2)||(sp3==2 && sp4==2 && sp5==2)||( sp6==2 && sp7==2 && sp8==2)||(sp0==2 && sp3==2 && sp6==2)||
    (sp1==2 && sp4==2 && sp7==2)||(sp2==2 && sp5==2 && sp8==2)||(sp0==2 && sp4==2 && sp8==2)||(sp2==2 && sp4==2 && sp6==2))
        win=2'b10;
    else if(sp0!=0 && sp1!=0 && sp2!=0 && sp3!=0 && sp4!=0 && sp5!=0 && sp6!=0 && sp7!=0 && sp8!=0)
        win=2'b11;
    else
        win=0;
end
end
endmodule

// GAME FSM
module game_fsm(sys_clk,reset,up,dn,rt,lt,select_x,select_y,enter,sp0,sp1,sp2,sp3,sp4,sp5,sp6,sp7,sp8,win);
input sys_clk,reset,up,dn,lt,rt,enter;
input [1:0]win;
output reg [9:0]select_x,select_y;
parameter s0=0,s1=1,s2=2,s3=3,s4=4,s5=5,s6=6,s7=7,s8=8;
parameter   box_h1=379,
            box_v1=108,
            box_h2=510,
            box_h3=640,
            box_v2=238,
            box_v3=368
            ;
reg [3:0]ps=s4;
reg [3:0]ns;
reg stop;
output reg [1:0]sp0=0,sp1=0,sp2=0,sp3=0,sp4=0,sp5=0,sp6=0,sp7=0,sp8=0;
always@(posedge sys_clk)
begin
if(reset)
begin
    ps<=s4;
end
else
begin 
    ps<=ns;
end
end
always@(posedge sys_clk)
begin
case(ps)
s0:if(up)
    ns<=s6;
    else if(lt)
    ns<=s2;
    else if(rt)
    ns<=s1;
    else if(dn)
    ns<=s3;
s1:if(up)
    ns<=s7;
    else if(lt)
    ns<=s0;
    else if(rt)
    ns<=s2;
    else if(dn)
    ns<=s4;
s2:if(up)
    ns<=s8;
    else if(lt)
    ns<=s1;
    else if(rt)
    ns<=s0;
    else if(dn)
    ns<=s5;
s3:if(up)
    ns<=s0;
    else if(lt)
    ns<=s5;
    else if(rt)
    ns<=s4;
    else if(dn)
    ns<=s6;
s4:if(up)
    ns<=s1;
    else if(lt)
    ns<=s3;
    else if(rt)
    ns<=s5;
    else if(dn)
    ns<=s7;
s5:if(up)
    ns<=s2;
    else if(lt)
    ns<=s4;
    else if(rt)
    ns<=s3;
    else if(dn)
    ns<=s8;
s6:if(up)
    ns<=s3;
    else if(lt)
    ns<=s8;
    else if(rt)
    ns<=s7;
    else if(dn)
    ns<=s0;
s7:if(up)
    ns<=s4;
    else if(lt)
    ns<=s6;
    else if(rt)
    ns<=s8;
    else if(dn)
    ns<=s1;
s8:if(up)
    ns<=s5;
    else if(lt)
    ns<=s7;
    else if(rt)
    ns<=s6;
    else if(dn)
    ns<=s2;
default:ns<=s4;
endcase
end
always@(posedge sys_clk)
begin
case(ps)
s0:begin 
   select_x=box_h1;
   select_y=box_v1;
   end 
s1:begin 
   select_x=box_h2;
   select_y=box_v1;
   end
s2:begin 
   select_x=box_h3;
   select_y=box_v1;
   end
s3:begin 
   select_x=box_h1;
   select_y=box_v2;
   end 
s4:begin 
   select_x=box_h2;
   select_y=box_v2;
   end
s5:begin 
   select_x=box_h3;
   select_y=box_v2;
   end
s6:begin 
   select_x=box_h1;
   select_y=box_v3;
   end 
s7:begin 
   select_x=box_h2;
   select_y=box_v3;
   end
s8:begin 
   select_x=box_h3;
   select_y=box_v3;
   end
default:
begin
    select_x=box_h1;
    select_y=box_v1;
end
endcase
end
reg person=1;
always@(posedge sys_clk)
begin
if(reset)
begin
    sp0=0;
    sp1=0;
    sp2=0;
    sp3=0;
    sp4=0;
    sp5=0;
    sp6=0;
    sp7=0;
    sp8=0;
    stop<=0;
    person<=1;
end
else
begin
    if(win>=1)
    stop=1;
    case(ps)
    s0:if(enter && sp0==0 && ~stop)
        begin
        person=person+1;
        if(person==0)
            sp0=1;
        else
            sp0=2;
        end
        else
        sp0=sp0;
    s1:if(enter && sp1==0 && ~stop)
        begin
        person=person+1;
        if(person==0)
            sp1=1;
        else
            sp1=2;
        end
        else
        sp1=sp1;
    s2:if(enter && sp2==0 && ~stop)
        begin
        person=person+1;
        if(person==0)
            sp2=1;
        else
            sp2=2;
        end
        else
        sp2=sp2;
    s3:if(enter && sp3==0 && ~stop)
        begin
        person=person+1;
        if(person==0)
            sp3=1;
        else
            sp3=2;
        end
        else
        sp3=sp3;
    s4:if(enter && sp4==0 && ~stop)
        begin
        person=person+1;
        if(person==0)
            sp4=1;
        else
            sp4=2;
        end
        else
        sp4=sp4;
    s5:if(enter && sp5==0 && ~stop)
        begin
        person=person+1;
        if(person==0)
            sp5=1;
        else
            sp5=2;
        end
        else
        sp5=sp5;
    s6:if(enter && sp6==0 && ~stop)
        begin
        person=person+1;
        if(person==0)
            sp6=1;
        else
            sp6=2;
        end
        else
        sp6=sp6;
    s7:if(enter && sp7==0 && ~stop)
        begin
        person=person+1;
        if(person==0)
            sp7=1;
        else
            sp7=2;
        end
        else
        sp7=sp7;
    s8:if(enter && sp8==0 && ~stop)
        begin
        person=person+1;
        if(person==0)
            sp8=1;
        else
            sp8=2;
        end
        else
        sp8=sp8;
    endcase
end
end 
endmodule

module DATA_TTT(clk_25M,data,head_adrs,data_sel);
input [6:0] head_adrs;
input clk_25M;
input [1:0]data_sel;
output reg [0:119]data;
always @(posedge clk_25M)
begin
case(data_sel)
1:case(head_adrs)
        7'd01:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd02:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd03:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd04:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd05:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd06:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd07:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd08:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd09:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd10:data<=100'b0000000000000000000111111111111111111000000000000000000000000000000000000011111111111111111000000000000000;
        7'd11:data<=100'b0000000000000000001111111111111111111100000000000000000000000000000000000111111111111111111100000000000000;
        7'd12:data<=100'b0000000000000000011111111111111111111110000000000000000000000000000000001111111111111111111100000000000000;
        7'd13:data<=100'b0000000000000000001111111111111111111110000000000000000000000000000000001111111111111111111100000000000000;
        7'd14:data<=100'b0000000000000000001111111111111111111111000000000000000000000000000000011111111111111111111100000000000000;
        7'd15:data<=100'b0000000000000000001111111111111111111111000000000000000000000000000000011111111111111111111000000000000000;
        7'd16:data<=100'b0000000000000000000111111111111111111111100000000000000000000000000000111111111111111111111000000000000000;
        7'd17:data<=100'b0000000000000000000111111111111111111111100000000000000000000000000000111111111111111111110000000000000000;
        7'd18:data<=100'b0000000000000000000011111111111111111111110000000000000000000000000001111111111111111111110000000000000000;
        7'd19:data<=100'b0000000000000000000001111111111111111111111000000000000000000000000001111111111111111111100000000000000000;
        7'd20:data<=100'b0000000000000000000001111111111111111111111000000000000000000000000011111111111111111111100000000000000000;
        7'd21:data<=100'b0000000000000000000000111111111111111111111100000000000000000000000011111111111111111111000000000000000000;
        7'd22:data<=100'b0000000000000000000000111111111111111111111100000000000000000000000111111111111111111111000000000000000000;
        7'd23:data<=100'b0000000000000000000000011111111111111111111110000000000000000000001111111111111111111110000000000000000000;
        7'd24:data<=100'b0000000000000000000000011111111111111111111110000000000000000000001111111111111111111100000000000000000000;
        7'd25:data<=100'b0000000000000000000000001111111111111111111111000000000000000000011111111111111111111100000000000000000000;
        7'd26:data<=100'b0000000000000000000000001111111111111111111111000000000000000000011111111111111111111000000000000000000000;
        7'd27:data<=100'b0000000000000000000000000111111111111111111111100000000000000000111111111111111111111000000000000000000000;
        7'd28:data<=100'b0000000000000000000000000111111111111111111111100000000000000000111111111111111111110000000000000000000000;
        7'd29:data<=100'b0000000000000000000000000011111111111111111111110000000000000001111111111111111111110000000000000000000000;
        7'd30:data<=100'b0000000000000000000000000001111111111111111111110000000000000001111111111111111111100000000000000000000000;
        7'd31:data<=100'b0000000000000000000000000001111111111111111111111000000000000011111111111111111111100000000000000000000000;
        7'd32:data<=100'b0000000000000000000000000000111111111111111111111000000000000011111111111111111111000000000000000000000000;
        7'd33:data<=100'b0000000000000000000000000000111111111111111111111100000000000111111111111111111110000000000000000000000000;
        7'd34:data<=100'b0000000000000000000000000000011111111111111111111110000000000111111111111111111110000000000000000000000000;
        7'd35:data<=100'b0000000000000000000000000000011111111111111111111110000000001111111111111111111100000000000000000000000000;
        7'd36:data<=100'b0000000000000000000000000000001111111111111111111111000000001111111111111111111100000000000000000000000000;
        7'd37:data<=100'b0000000000000000000000000000001111111111111111111111000000011111111111111111111000000000000000000000000000;
        7'd38:data<=100'b0000000000000000000000000000000111111111111111111111100000011111111111111111111000000000000000000000000000;
        7'd39:data<=100'b0000000000000000000000000000000111111111111111111111100000111111111111111111110000000000000000000000000000;
        7'd40:data<=100'b0000000000000000000000000000000011111111111111111111110000111111111111111111110000000000000000000000000000;
        7'd41:data<=100'b0000000000000000000000000000000001111111111111111111110001111111111111111111100000000000000000000000000000;
        7'd42:data<=100'b0000000000000000000000000000000001111111111111111111111001111111111111111111100000000000000000000000000000;
        7'd43:data<=100'b0000000000000000000000000000000000111111111111111111111011111111111111111111000000000000000000000000000000;
        7'd44:data<=100'b0000000000000000000000000000000000111111111111111111111111111111111111111110000000000000000000000000000000;
        7'd45:data<=100'b0000000000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000;
        7'd46:data<=100'b0000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000000000000000;
        7'd47:data<=100'b0000000000000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000;
        7'd48:data<=100'b0000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000000000000;
        7'd49:data<=100'b0000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000000000000000000;
        7'd50:data<=100'b0000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000000;
        7'd51:data<=100'b0000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000000000000000000;
        7'd52:data<=100'b0000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000;
        7'd53:data<=100'b0000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000;
        7'd54:data<=100'b0000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000;
        7'd55:data<=100'b0000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000;
        7'd56:data<=100'b0000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000;
        7'd57:data<=100'b0000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000;
        7'd58:data<=100'b0000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000;
        7'd59:data<=100'b0000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000;
        7'd60:data<=100'b0000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000;
        7'd61:data<=100'b0000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000;
        7'd62:data<=100'b0000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000000000000000000;
        7'd63:data<=100'b0000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000000;
        7'd64:data<=100'b0000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000000000000000000;
        7'd65:data<=100'b0000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000000000000;
        7'd66:data<=100'b0000000000000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000;
        7'd67:data<=100'b0000000000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000;
        7'd68:data<=100'b0000000000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000;
        7'd69:data<=100'b0000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000;
        7'd70:data<=100'b0000000000000000000000000000000000111111111111111111110111111111111111111111000000000000000000000000000000;
        7'd71:data<=100'b0000000000000000000000000000000001111111111111111111100111111111111111111111100000000000000000000000000000;
        7'd72:data<=100'b0000000000000000000000000000000011111111111111111111100011111111111111111111100000000000000000000000000000;
        7'd73:data<=100'b0000000000000000000000000000000011111111111111111111000011111111111111111111110000000000000000000000000000;
        7'd74:data<=100'b0000000000000000000000000000000111111111111111111110000001111111111111111111110000000000000000000000000000;
        7'd75:data<=100'b0000000000000000000000000000000111111111111111111110000001111111111111111111111000000000000000000000000000;
        7'd76:data<=100'b0000000000000000000000000000001111111111111111111100000000111111111111111111111000000000000000000000000000;
        7'd77:data<=100'b0000000000000000000000000000001111111111111111111100000000111111111111111111111100000000000000000000000000;
        7'd78:data<=100'b0000000000000000000000000000011111111111111111111000000000011111111111111111111100000000000000000000000000;
        7'd79:data<=100'b0000000000000000000000000000011111111111111111111000000000011111111111111111111110000000000000000000000000;
        7'd80:data<=100'b0000000000000000000000000000111111111111111111110000000000001111111111111111111111000000000000000000000000;
        7'd81:data<=100'b0000000000000000000000000001111111111111111111110000000000001111111111111111111111000000000000000000000000;
        7'd82:data<=100'b0000000000000000000000000001111111111111111111100000000000000111111111111111111111100000000000000000000000;
        7'd83:data<=100'b0000000000000000000000000011111111111111111111100000000000000111111111111111111111100000000000000000000000;
        7'd84:data<=100'b0000000000000000000000000011111111111111111111000000000000000011111111111111111111110000000000000000000000;
        7'd85:data<=100'b0000000000000000000000000111111111111111111111000000000000000001111111111111111111110000000000000000000000;
        7'd86:data<=100'b0000000000000000000000000111111111111111111110000000000000000001111111111111111111111000000000000000000000;
        7'd87:data<=100'b0000000000000000000000001111111111111111111110000000000000000000111111111111111111111000000000000000000000;
        7'd88:data<=100'b0000000000000000000000001111111111111111111100000000000000000000111111111111111111111100000000000000000000;
        7'd89:data<=100'b0000000000000000000000011111111111111111111100000000000000000000011111111111111111111100000000000000000000;
        7'd90:data<=100'b0000000000000000000000011111111111111111111000000000000000000000011111111111111111111110000000000000000000;
        7'd91:data<=100'b0000000000000000000000111111111111111111111000000000000000000000001111111111111111111111000000000000000000;
        7'd92:data<=100'b0000000000000000000001111111111111111111110000000000000000000000001111111111111111111111000000000000000000;
        7'd93:data<=100'b0000000000000000000001111111111111111111110000000000000000000000000111111111111111111111100000000000000000;
        7'd94:data<=100'b0000000000000000000011111111111111111111100000000000000000000000000111111111111111111111100000000000000000;
        7'd95:data<=100'b0000000000000000000011111111111111111111100000000000000000000000000011111111111111111111110000000000000000;
        7'd96:data<=100'b0000000000000000000111111111111111111111000000000000000000000000000011111111111111111111110000000000000000;
        7'd97:data<=100'b0000000000000000000111111111111111111110000000000000000000000000000001111111111111111111111000000000000000;
        7'd98:data<=100'b0000000000000000001111111111111111111110000000000000000000000000000001111111111111111111111000000000000000;
        7'd99:data<=100'b0000000000000000001111111111111111111100000000000000000000000000000000111111111111111111111100000000000000;
        7'd100:data<=100'b0000000000000000011111111111111111111100000000000000000000000000000000111111111111111111111100000000000000;
        7'd101:data<=100'b0000000000000000011111111111111111111000000000000000000000000000000000011111111111111111111110000000000000;
        7'd102:data<=100'b0000000000000000111111111111111111111000000000000000000000000000000000011111111111111111111110000000000000;
        7'd103:data<=100'b0000000000000000111111111111111111110000000000000000000000000000000000001111111111111111111110000000000000;
        7'd104:data<=100'b0000000000000000111111111111111111110000000000000000000000000000000000001111111111111111111110000000000000;
        7'd105:data<=100'b0000000000000000111111111111111111100000000000000000000000000000000000000111111111111111111110000000000000;
        7'd106:data<=100'b00000000000000001111111111111111111000000000000000000000000000000000000000111111111111111110000000000000000;
        7'd107:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd108:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd109:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd110:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd111:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd112:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd113:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


    endcase
2:case(head_adrs)
        7'd01:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd02:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd03:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd04:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd05:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd06:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd07:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd08:data<=100'b00000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000;
        7'd09:data<=100'b00000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000;
        7'd10:data<=100'b00000000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000000000000000;
        7'd11:data<=100'b00000000000000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000;
        7'd12:data<=100'b00000000000000000000000000000000000001111111111111111111111111111111111111111111110000000000000000000000000;
        7'd13:data<=100'b00000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000;
        7'd14:data<=100'b00000000000000000000000000000000011111111111111111111111111111111111111111111111111110000000000000000000000;
        7'd15:data<=100'b00000000000000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000;
        7'd16:data<=100'b00000000000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000000000000;
        7'd17:data<=100'b00000000000000000000000000000111111111111111111111111111111111111111111111111111111111111100000000000000000;
        7'd18:data<=100'b00000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000;
        7'd19:data<=100'b00000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000;
        7'd20:data<=100'b00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000;
        7'd21:data<=100'b00000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000;
        7'd22:data<=100'b00000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000;
        7'd23:data<=100'b00000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111000000000000;
        7'd24:data<=100'b00000000000000000000001111111111111111111111111111111110000001111111111111111111111111111111111100000000000;
        7'd25:data<=100'b00000000000000000000011111111111111111111111111111000000000000000001111111111111111111111111111100000000000;
        7'd26:data<=100'b00000000000000000000111111111111111111111111111000000000000000000000011111111111111111111111111110000000000;
        7'd27:data<=100'b00000000000000000000111111111111111111111111100000000000000000000000000111111111111111111111111111000000000;
        7'd28:data<=100'b00000000000000000001111111111111111111111111000000000000000000000000000001111111111111111111111111000000000;
        7'd29:data<=100'b00000000000000000011111111111111111111111110000000000000000000000000000000111111111111111111111111100000000;
        7'd30:data<=100'b00000000000000000011111111111111111111111000000000000000000000000000000000011111111111111111111111100000000;
        7'd31:data<=100'b00000000000000000111111111111111111111110000000000000000000000000000000000001111111111111111111111100000000;
        7'd32:data<=100'b00000000000000000111111111111111111111110000000000000000000000000000000000000111111111111111111111110000000;
        7'd33:data<=100'b00000000000000000111111111111111111111100000000000000000000000000000000000000011111111111111111111110000000;
        7'd34:data<=100'b00000000000000001111111111111111111111000000000000000000000000000000000000000011111111111111111111111000000;
        7'd35:data<=100'b00000000000000001111111111111111111110000000000000000000000000000000000000000001111111111111111111111000000;
        7'd36:data<=100'b00000000000000011111111111111111111110000000000000000000000000000000000000000001111111111111111111111000000;
        7'd37:data<=100'b00000000000000011111111111111111111100000000000000000000000000000000000000000000111111111111111111111100000;
        7'd38:data<=100'b00000000000000011111111111111111111100000000000000000000000000000000000000000000111111111111111111111100000;
        7'd39:data<=100'b00000000000000111111111111111111111100000000000000000000000000000000000000000000011111111111111111111100000;
        7'd40:data<=100'b00000000000000111111111111111111111000000000000000000000000000000000000000000000011111111111111111111100000;
        7'd41:data<=100'b00000000000000111111111111111111111000000000000000000000000000000000000000000000011111111111111111111100000;
        7'd42:data<=100'b00000000000000111111111111111111111000000000000000000000000000000000000000000000011111111111111111111110000;
        7'd43:data<=100'b00000000000001111111111111111111110000000000000000000000000000000000000000000000001111111111111111111110000;
        7'd44:data<=100'b00000000000001111111111111111111110000000000000000000000000000000000000000000000001111111111111111111110000;
        7'd45:data<=100'b00000000000001111111111111111111110000000000000000000000000000000000000000000000001111111111111111111110000;
        7'd46:data<=100'b00000000000001111111111111111111110000000000000000000000000000000000000000000000001111111111111111111110000;
        7'd47:data<=100'b00000000000001111111111111111111100000000000000000000000000000000000000000000000001111111111111111111110000;
        7'd48:data<=100'b00000000000001111111111111111111100000000000000000000000000000000000000000000000000111111111111111111110000;
        7'd49:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111110000;
        7'd50:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd51:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd52:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd53:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd54:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd55:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd56:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd57:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd58:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd59:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd60:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd61:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd62:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd63:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd64:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111000;
        7'd65:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111110000;
        7'd66:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111110000;
        7'd67:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000000111111111111111111110000;
        7'd68:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000001111111111111111111110000;
        7'd69:data<=100'b00000000000011111111111111111111100000000000000000000000000000000000000000000000001111111111111111111110000;
        7'd70:data<=100'b00000000000001111111111111111111100000000000000000000000000000000000000000000000001111111111111111111110000;
        7'd71:data<=100'b00000000000001111111111111111111110000000000000000000000000000000000000000000000001111111111111111111110000;
        7'd72:data<=100'b00000000000001111111111111111111110000000000000000000000000000000000000000000000001111111111111111111110000;
        7'd73:data<=100'b00000000000001111111111111111111110000000000000000000000000000000000000000000000001111111111111111111100000;
        7'd74:data<=100'b00000000000001111111111111111111110000000000000000000000000000000000000000000000011111111111111111111100000;
        7'd75:data<=100'b00000000000001111111111111111111110000000000000000000000000000000000000000000000011111111111111111111100000;
        7'd76:data<=100'b00000000000001111111111111111111111000000000000000000000000000000000000000000000011111111111111111111100000;
        7'd77:data<=100'b00000000000000111111111111111111111000000000000000000000000000000000000000000000111111111111111111111000000;
        7'd78:data<=100'b00000000000000111111111111111111111000000000000000000000000000000000000000000000111111111111111111111000000;
        7'd79:data<=100'b00000000000000111111111111111111111100000000000000000000000000000000000000000000111111111111111111111000000;
        7'd80:data<=100'b00000000000000111111111111111111111100000000000000000000000000000000000000000001111111111111111111110000000;
        7'd81:data<=100'b00000000000000011111111111111111111110000000000000000000000000000000000000000001111111111111111111110000000;
        7'd82:data<=100'b00000000000000011111111111111111111110000000000000000000000000000000000000000011111111111111111111110000000;
        7'd83:data<=100'b00000000000000011111111111111111111111000000000000000000000000000000000000000111111111111111111111100000000;
        7'd84:data<=100'b00000000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111100000000;
        7'd85:data<=100'b00000000000000001111111111111111111111100000000000000000000000000000000000001111111111111111111111100000000;
        7'd86:data<=100'b00000000000000001111111111111111111111110000000000000000000000000000000000011111111111111111111111000000000;
        7'd87:data<=100'b00000000000000000111111111111111111111111000000000000000000000000000000000111111111111111111111111000000000;
        7'd88:data<=100'b00000000000000000111111111111111111111111100000000000000000000000000000001111111111111111111111110000000000;
        7'd89:data<=100'b00000000000000000011111111111111111111111110000000000000000000000000000111111111111111111111111100000000000;
        7'd90:data<=100'b00000000000000000011111111111111111111111111100000000000000000000000001111111111111111111111111100000000000;
        7'd91:data<=100'b00000000000000000001111111111111111111111111111000000000000000000001111111111111111111111111111000000000000;
        7'd92:data<=100'b00000000000000000001111111111111111111111111111111100000000000001111111111111111111111111111110000000000000;
        7'd93:data<=100'b00000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111110000000000000;
        7'd94:data<=100'b00000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000;
        7'd95:data<=100'b00000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111000000000000000;
        7'd96:data<=100'b00000000000000000000001111111111111111111111111111111111111111111111111111111111111111111110000000000000000;
        7'd97:data<=100'b00000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000000000000;
        7'd98:data<=100'b00000000000000000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000;
        7'd99:data<=100'b00000000000000000000000001111111111111111111111111111111111111111111111111111111111111110000000000000000000;
        7'd100:data<=100'b00000000000000000000000000011111111111111111111111111111111111111111111111111111111111100000000000000000000;
        7'd101:data<=100'b00000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000;
        7'd102:data<=100'b00000000000000000000000000000111111111111111111111111111111111111111111111111111111100000000000000000000000;
        7'd103:data<=100'b00000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000;
        7'd104:data<=100'b00000000000000000000000000000000011111111111111111111111111111111111111111111111000000000000000000000000000;
        7'd105:data<=100'b00000000000000000000000000000000000111111111111111111111111111111111111111111100000000000000000000000000000;
        7'd106:data<=100'b00000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000;
        7'd107:data<=100'b00000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000000000000;
        7'd108:data<=100'b00000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000;
        7'd109:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd110:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd111:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd112:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd113:data<=100'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
 default:case(head_adrs)
        7'd01:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd02:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd03:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd04:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd05:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd06:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd07:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd08:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd09:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd10:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd11:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd12:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd13:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd14:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd15:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd16:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd17:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd18:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd19:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd20:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd21:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd22:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd23:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd24:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd25:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd26:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd27:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd28:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd29:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd30:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd31:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd32:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd33:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd34:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd35:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd36:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd37:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd38:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd39:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd40:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd41:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd42:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd43:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd44:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd45:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd46:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd47:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd48:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd49:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd50:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd51:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd52:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd53:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd54:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd55:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd56:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd57:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd58:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd59:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd60:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd61:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd62:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd63:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd64:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd65:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd66:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd67:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd68:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd69:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd70:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd71:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd72:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd73:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd74:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd75:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd76:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd77:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd78:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd79:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd80:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd81:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd82:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd83:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd84:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd85:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd86:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd87:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd88:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd89:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd90:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd91:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd92:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd93:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd94:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd95:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd96:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd97:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd98:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd99:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd100:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd101:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd102:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd103:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd104:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd105:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd106:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd107:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd108:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd109:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd110:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd111:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd112:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7'd113:data<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
   endcase                              
 endcase
end
endmodule
module Title_TTT(clk_25M,title,title_adrs,player,player_adrs);
input clk_25M;
output reg [0:423] title;
input [6:0] player_adrs;
output reg [0:219] player;
input [5:0] title_adrs;
always @(posedge clk_25M)
begin
    case(title_adrs)
        6'd00:title<=424'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd01:title<=424'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000;
        6'd02:title<=424'b001111111111111111111111111111111111111100000001111111111000000000000000000000000001111111111111111100000000000000000000000000000000000111111111111111111111111111111111111100000000000000001111111111100000000000000000000000000000000000001111111111111111100000000000000000000000000000000001111111111111111111111111111111111111100000000000000000011111111111111111100000000000000000000000000111111111111111111111111111111111100;
        6'd03:title<=424'b001111111111111111111111111111111111111100000001111111111000000000000000000000000111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111100000000000000011111111111100000000000000000000000000000000001111111111111111111111100000000000000000000000000000001111111111111111111111111111111111111100000000000000001111111111111111111111100000000000000000000000111111111111111111111111111111111100;
        6'd04:title<=424'b001111111111111111111111111111111111111100000001111111111000000000000000000000011111111111111111111111111000000000000000000000000000000111111111111111111111111111111111111100000000000000011111111111110000000000000000000000000000000111111111111111111111111111000000000000000000000000000001111111111111111111111111111111111111100000000000000111111111111111111111111111000000000000000000000111111111111111111111111111111111100;
        6'd05:title<=424'b001111111111111111111111111111111111111100000001111111111000000000000000000001111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111100000000000000111111111111110000000000000000000000000000001111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111100000000000011111111111111111111111111111100000000000000000000111111111111111111111111111111111100;
        6'd06:title<=424'b001111111111111111111111111111111111111100000001111111111000000000000000000011111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111100000000000000111111111111111000000000000000000000000000111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111100000000000111111111111111111111111111111111000000000000000000111111111111111111111111111111111100;
        6'd07:title<=424'b001111111111111111111111111111111111111100000001111111111000000000000000000111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111100000000000000111111111111111000000000000000000000000001111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111100000000001111111111111111111111111111111111100000000000000000111111111111111111111111111111111100;
        6'd08:title<=424'b001111111111111111111111111111111111111100000001111111111000000000000000001111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111100000000000001111111111111111000000000000000000000000011111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111100000000011111111111111111111111111111111111110000000000000000111111111111111111111111111111111100;
        6'd09:title<=424'b001111111111111111111111111111111111111100000001111111111000000000000000011111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111100000000000001111111111111111100000000000000000000000111111111111111111111111111111111111111000000000000000000000001111111111111111111111111111111111111100000000111111111111111111111111111111111111111000000000000000111111111111111111111111111111111100;
        6'd10:title<=424'b001111111111111111111111111111111111111100000001111111111000000000000000111111111111111110000001111111111111111100000000000000000000000111111111111111111111111111111111111100000000000001111111111111111100000000000000000000000111111111111111100000001111111111111111000000000000000000000001111111111111111111111111111111111111100000001111111111111111100000001111111111111111000000000000000111111111111111111111111111111111100;
        6'd11:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000001111111111111110000000000001111111111111100000000000000000000000000000000000011111111111000000000000000000000000011111111111111111100000000000000000000001111111111111100000000000001111111111111100000000000000000000000000000000000011111111110000000000000000000001111111111111100000000000001111111111111100000000000000111111111110000000000000000000000000;
        6'd12:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000001111111111111000000000000000011111111111110000000000000000000000000000000000011111111111000000000000000000000000011111111111111111110000000000000000000011111111111110000000000000000111111111111100000000000000000000000000000000000011111111110000000000000000000011111111111110000000000000000111111111111110000000000000111111111110000000000000000000000000;
        6'd13:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000011111111111110000000000000000001111111111110000000000000000000000000000000000011111111111000000000000000000000000011111111111111111110000000000000000000011111111111100000000000000000011111111111110000000000000000000000000000000000011111111110000000000000000000011111111111100000000000000000011111111111110000000000000111111111110000000000000000000000000;
        6'd14:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000011111111111100000000000000000000111111111111000000000000000000000000000000000011111111111000000000000000000000000111111111101111111110000000000000000000111111111111000000000000000000001111111111110000000000000000000000000000000000011111111110000000000000000000111111111111000000000000000000001111111111111000000000000111111111110000000000000000000000000;
        6'd15:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000111111111111000000000000000000000111111111111000000000000000000000000000000000011111111111000000000000000000000000111111111001111111111000000000000000000111111111111000000000000000000000111111111110000000000000000000000000000000000011111111110000000000000000000111111111111000000000000000000000111111111111000000000000111111111110000000000000000000000000;
        6'd16:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000111111111111000000000000000000000011111111111000000000000000000000000000000000011111111111000000000000000000000001111111111000111111111000000000000000001111111111110000000000000000000000111111111111000000000000000000000000000000000011111111110000000000000000001111111111110000000000000000000000011111111111000000000000111111111110000000000000000000000000;
        6'd17:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000111111111110000000000000000000000011111111111000000000000000000000000000000000011111111111000000000000000000000001111111111000111111111000000000000000001111111111110000000000000000000000011111111111000000000000000000000000000000000011111111110000000000000000001111111111100000000000000000000000011111111111100000000000111111111110000000000000000000000000;
        6'd18:title<=424'b000000000000000011111111110000000000000000000001111111111000000000001111111111110000000000000000000000011111111111000000000000000000000000000000000011111111111000000000000000000000001111111110000111111111100000000000000001111111111100000000000000000000000011111111111000000000000000000000000000000000011111111110000000000000000001111111111100000000000000000000000001111111111100000000000111111111110000000000000000000000000;
        6'd19:title<=424'b000000000000000011111111110000000000000000000001111111111000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000011111111110000011111111100000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111100000000000000000000000001111111111100000000000111111111110000000000000000000000000;
        6'd20:title<=424'b000000000000000011111111110000000000000000000001111111111000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000011111111110000011111111110000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000001111111111100000000000111111111110000000000000000000000000;
        6'd21:title<=424'b000000000000000011111111110000000000000000000001111111111000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000011111111100000011111111110000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111110000000000000000000000000;
        6'd22:title<=424'b000000000000000011111111110000000000000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000111111111100000001111111110000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111110000000000000000000000000;
        6'd23:title<=424'b000000000000000011111111110000000000000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000111111111100000001111111111000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111111111111111111111111110000;
        6'd24:title<=424'b000000000000000011111111110000000000000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000111111111000000001111111111000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111111111111111111111111110000;
        6'd25:title<=424'b000000000000000011111111110000000000000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000001111111111000000000111111111000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111111111111111111111111110000;
        6'd26:title<=424'b000000000000000011111111110000000000000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000001111111111000000000111111111100000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111111111111111111111111110000;
        6'd27:title<=424'b000000000000000011111111110000000000000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000001111111110000000000111111111100000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111111111111111111111111110000;
        6'd28:title<=424'b000000000000000011111111110000000000000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000011111111110000000000111111111100000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111111111111111111111111110000;
        6'd29:title<=424'b000000000000000011111111110000000000000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000011111111110000000000011111111110000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111111111111111111111111110000;
        6'd30:title<=424'b000000000000000011111111110000000000000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000111111111100000000000011111111110000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111111111111111111111111110000;
        6'd31:title<=424'b000000000000000011111111110000000000000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000111111111100000000000011111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111110000000000000000000000000;
        6'd32:title<=424'b000000000000000011111111110000000000000000000001111111111000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000111111111100000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000000111111111110000000000111111111110000000000000000000000000;
        6'd33:title<=424'b000000000000000011111111110000000000000000000001111111111000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000001111111111111111111111111111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000001111111111110000000000111111111110000000000000000000000000;
        6'd34:title<=424'b000000000000000011111111110000000000000000000001111111111000000000001111111111100000000000000000000000001111111111000000000000000000000000000000000011111111111000000000000000001111111111111111111111111111111111100000000011111111111000000000000000000000000011111111111000000000000000000000000000000000011111111110000000000000000011111111111000000000000000000000000001111111111100000000000111111111110000000000000000000000000;
        6'd35:title<=424'b000000000000000011111111110000000000000000000001111111111000000000001111111111100000000000000000000000011111111111000000000000000000000000000000000011111111111000000000000000001111111111111111111111111111111111100000000011111111111100000000000000000000000011111111111000000000000000000000000000000000011111111110000000000000000011111111111100000000000000000000000001111111111100000000000111111111110000000000000000000000000;
        6'd36:title<=424'b000000000000000011111111110000000000000000000001111111111000000000001111111111110000000000000000000000011111111111000000000000000000000000000000000011111111111000000000000000011111111111111111111111111111111111100000000001111111111100000000000000000000000011111111111000000000000000000000000000000000011111111110000000000000000001111111111100000000000000000000000001111111111100000000000111111111110000000000000000000000000;
        6'd37:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000111111111110000000000000000000000011111111111000000000000000000000000000000000011111111111000000000000000011111111111111111111111111111111111110000000001111111111110000000000000000000000011111111111000000000000000000000000000000000011111111110000000000000000001111111111100000000000000000000000011111111111100000000000111111111110000000000000000000000000;
        6'd38:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000111111111111000000000000000000000011111111111000000000000000000000000000000000011111111111000000000000000011111111111111111111111111111111111110000000001111111111110000000000000000000000111111111110000000000000000000000000000000000011111111110000000000000000001111111111110000000000000000000000011111111111000000000000111111111110000000000000000000000000;
        6'd39:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000111111111111000000000000000000000111111111111000000000000000000000000000000000011111111111000000000000000111111111111111111111111111111111111110000000000111111111111000000000000000000000111111111110000000000000000000000000000000000011111111110000000000000000000111111111111000000000000000000000111111111111000000000000111111111110000000000000000000000000;
        6'd40:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000011111111111100000000000000000001111111111110000000000000000000000000000000000011111111111000000000000000111111111111111111111111111111111111111000000000111111111111000000000000000000001111111111110000000000000000000000000000000000011111111110000000000000000000111111111111000000000000000000001111111111111000000000000111111111110000000000000000000000000;
        6'd41:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000011111111111110000000000000000001111111111110000000000000000000000000000000000011111111111000000000000000111111111111111111111111111111111111111000000000011111111111100000000000000000011111111111100000000000000000000000000000000000011111111110000000000000000000011111111111100000000000000000011111111111110000000000000111111111110000000000000000000000000;
        6'd42:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000001111111111111000000000000000111111111111110000000000000000000000000000000000011111111111000000000000001111111111100000000000000000001111111111000000000011111111111111000000000000000111111111111100000000000000000000000000000000000011111111110000000000000000000011111111111111000000000000000111111111111110000000000000111111111110000000000000000000000000;
        6'd43:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000001111111111111110000000000001111111111111100000000000000000000000000000000000011111111111000000000000001111111111100000000000000000001111111111100000000001111111111111100000000000011111111111111100000000000000000000000000000000000011111111110000000000000000000001111111111111100000000000011111111111111100000000000000111111111110000000000000000000000000;
        6'd44:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000000111111111111111110000011111111111111111000000000000000000000000000000000000011111111111000000000000011111111111000000000000000000001111111111100000000000111111111111111110000011111111111111111000000000000000000000000000000000000011111111110000000000000000000001111111111111111110000011111111111111111000000000000000111111111111111111111111111111111100;
        6'd45:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000011111111111000000000000011111111111000000000000000000000111111111110000000000111111111111111111111111111111111111110000000000000000000000000000000000000011111111110000000000000000000000111111111111111111111111111111111111110000000000000000111111111111111111111111111111111100;
        6'd46:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000000001111111111111111111111111111111111110000000000000000000000000000000000000011111111111000000000000011111111111000000000000000000000111111111110000000000011111111111111111111111111111111111110000000000000000000000000000000000000011111111110000000000000000000000011111111111111111111111111111111111110000000000000000111111111111111111111111111111111100;
        6'd47:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000000000111111111111111111111111111111111100000000000000000000000000000000000000011111111111000000000000111111111110000000000000000000000111111111110000000000001111111111111111111111111111111111100000000000000000000000000000000000000011111111110000000000000000000000001111111111111111111111111111111111100000000000000000111111111111111111111111111111111100;
        6'd48:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000011111111111000000000000111111111110000000000000000000000011111111111000000000000111111111111111111111111111111111000000000000000000000000000000000000000011111111110000000000000000000000000111111111111111111111111111111110000000000000000000111111111111111111111111111111111100;
        6'd49:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000011111111111000000000000111111111110000000000000000000000011111111111000000000000001111111111111111111111111111100000000000000000000000000000000000000000011111111110000000000000000000000000001111111111111111111111111111100000000000000000000111111111111111111111111111111111100;
        6'd50:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000011111111111000000000001111111111100000000000000000000000011111111111000000000000000111111111111111111111111111000000000000000000000000000000000000000000011111111110000000000000000000000000000111111111111111111111111111000000000000000000000111111111111111111111111111111111100;
        6'd51:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000011111111111000000000001111111111100000000000000000000000001111111111100000000000000001111111111111111111111100000000000000000000000000000000000000000000011111111110000000000000000000000000000001111111111111111111111100000000000000000000000111111111111111111111111111111111100;
        6'd52:title<=424'b000000000000000011111111110000000000000000000001111111111000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000011111111111000000000001111111111000000000000000000000000001111111111100000000000000000001111111111111111100000000000000000000000000000000000000000000000011111111110000000000000000000000000000000001111111111111111100000000000000000000000000111111111111111111111111111111111100;
        6'd53:title<=424'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000;
        6'd54:title<=424'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        default: title<=0;
    endcase
end
always @(posedge clk_25M)
begin
    case(player_adrs)
    7'd00:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd01:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd02:player<=220'b0111111111111100000000001111100000000000000000000011111100000001111110000000000111111000111111111111111110000011111111111111100000000000000000000000000000000000000000000000000000000000000000000011111100000000011111100000;
7'd03:player<=220'b0111111111111111000000001111100000000000000000000011111100000001111110000000000111110000111111111111111110000011111111111111110000000000000000000000011111000000000000000000000000000000000000000001111110000000011111000000;
7'd04:player<=220'b0111111111111111100000001111100000000000000000000111111110000000111111000000001111110000111111111111111110000011111111111111111000000000000000000000111111000000000000000000000000000000000000000001111110000000111111000000;
7'd05:player<=220'b0111111111111111110000001111100000000000000000000111111110000000111111000000001111110000111111111111111110000011111111111111111100000000000000000001111111000000000000000000000000000000000000000000111111000000111110000000;
7'd06:player<=220'b0111111111111111110000001111100000000000000000000111111110000000011111000000011111100000111111111111111110000011111111111111111100000000000000000011111111000000000000000000000000000000000000000000111111000001111110000000;
7'd07:player<=220'b0111110000011111111000001111100000000000000000000111111110000000011111100000011111100000111111000000000000000011111100000111111110000000000000001111111111000000000000000000000000000000000000000000011111000001111100000000;
7'd08:player<=220'b0111110000000111111000001111100000000000000000001111111111000000011111100000011111000000111110000000000000000011111000000001111110000000000000111111111111000000000000000000000000000000000000000000011111100011111100000000;
7'd09:player<=220'b0111110000000011111000001111100000000000000000001111111111000000001111100000111111000000111110000000000000000011111000000001111110000000000000111111111111000000000000000000000000000000000000000000001111100011111000000000;
7'd10:player<=220'b0111110000000011111000001111100000000000000000001111001111000000001111110000111110000000111110000000000000000011111000000000111110000000000000111111111111000000000000000000000000000000000000000000001111110111111000000000;
7'd11:player<=220'b0111110000000011111000001111100000000000000000001111001111100000000111110000111110000000111110000000000000000011111000000000111110000000000000111110011111000000000000000000000000000000000000000000000111110111110000000000;
7'd12:player<=220'b0111110000000011111100001111100000000000000000011111001111100000000111111001111110000000111110000000000000000011111000000000111110000000000000111100011111000000000000000000000000000000000000000000000111111111110000000000;
7'd13:player<=220'b0111110000000011111000001111100000000000000000011111001111100000000011111001111100000000111110000000000000000011111000000001111110000000000000110000011111000000000000000000000000000000000000000000000011111111100000000000;
7'd14:player<=220'b0111110000000011111000001111100000000000000000011110000111100000000011111011111100000000111111000000000000000011111000000001111100000000000000000000011111000000000000000000000000000000000000000000000011111111100000000000;
7'd15:player<=220'b0111110000000111111000001111100000000000000000111110000111110000000011111111111000000000111111111111111100000011111000000011111100000000000000000000011111000000000000000000000000000000000000000000000001111111000000000000;
7'd16:player<=220'b0111110000001111111000001111100000000000000000111110000111110000000001111111111000000000111111111111111100000011111111111111111000000000000000000000011111000000000000000000000000000000000000000000000001111111000000000000;
7'd17:player<=220'b0111111111111111111000001111100000000000000000111110000111110000000001111111111000000000111111111111111100000011111111111111110000000000000000000000011111000000000000000000000000000000000000000000000001111111000000000000;
7'd18:player<=220'b0111111111111111110000001111100000000000000000111100000011110000000000111111110000000000111111111111111100000011111111111111100000000000000000000000011111000000000000000000000000000000000000000000000001111111000000000000;
7'd19:player<=220'b0111111111111111100000001111100000000000000001111100000011111000000000111111110000000000111111111111111100000011111111111111100000000000000000000000011111000000000000000000000000000000000000000000000001111111100000000000;
7'd20:player<=220'b0111111111111111000000001111100000000000000001111100000011111000000000011111100000000000111111000000000000000011111111111111111000000000000000000000011111000000000000001111111111111111100000000000000011111111100000000000;
7'd21:player<=220'b0111111111111110000000001111100000000000000001111111111111111000000000011111100000000000111110000000000000000011111111111111111000000000000000000000011111000000000000001111111111111111100000000000000011111111110000000000;
7'd22:player<=220'b0111111111110000000000001111100000000000000011111111111111111100000000011111100000000000111110000000000000000011111000000011111100000000000000000000011111000000000000001111111111111111100000000000000111111111110000000000;
7'd23:player<=220'b0111110000000000000000001111100000000000000011111111111111111100000000011111100000000000111110000000000000000011111000000001111100000000000000000000011111000000000000001111111111111111100000000000000111111111111000000000;
7'd24:player<=220'b0111110000000000000000001111100000000000000011111111111111111100000000011111100000000000111110000000000000000011111000000001111110000000000000000000011111000000000000001111111111111111100000000000001111110111111000000000;
7'd25:player<=220'b0111110000000000000000001111100000000000000011111111111111111100000000011111100000000000111110000000000000000011111000000001111110000000000000000000011111000000000000000000000000000000000000000000001111100011111100000000;
7'd26:player<=220'b0111110000000000000000001111100000000000000111111111111111111110000000011111100000000000111110000000000000000011111000000000111110000000000000000000011111000000000000000000000000000000000000000000011111100011111100000000;
7'd27:player<=220'b0111110000000000000000001111100000000000000111110000000000111110000000011111100000000000111110000000000000000011111000000000111110000000000000000000011111000000000000000000000000000000000000000000011111000001111110000000;
7'd28:player<=220'b0111110000000000000000001111111111111111000111110000000000111110000000011111100000000000111111000000000000000011111000000000111110000000000000000000011111000000000000000000000000000000000000000000111111000001111110000000;
7'd29:player<=220'b0111110000000000000000001111111111111111000111110000000000111111000000011111100000000000111111111111111110000011111000000000111111000000000000000000011111000000000000000000000000000000000000000000111110000000111111000000;
7'd30:player<=220'b0111110000000000000000001111111111111111001111110000000000111111000000011111100000000000111111111111111110000011111000000000111111000000000000000000011111000000000000000000000000000000000000000001111110000000111111000000;
7'd31:player<=220'b0111110000000000000000001111111111111111001111100000000000011111000000011111100000000000111111111111111110000011111000000000011111000000000000000000011111000000000000000000000000000000000000000001111100000000111111100000;
7'd32:player<=220'b0111110000000000000000001111111111111111001111100000000000011111000000011111100000000000111111111111111110000011111000000000011111000000000000000000011111000000000000000000000000000000000000000011111100000000011111100000;
7'd33:player<=220'b0111110000000000000000001111111111111111011111100000000000011111100000011111100000000000111111111111111110000011111000000000011111100000000000000000011111000000000000000000000000000000000000000011111000000000011111110000;
7'd34:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd35:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd36:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd37:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd38:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd39:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd40:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd41:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd42:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd43:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd44:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd45:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd46:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd47:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd48:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000;
7'd49:player<=220'b0111111111111100000000001111100000000000000000000011111100000001111110000000000111111000111111111111111110000011111111111111000000000000000000000000111000000000000000000000000000000000000000000000000000111111111100000000;
7'd50:player<=220'b0111111111111111000000001111100000000000000000000011111100000001111110000000000111110000111111111111111110000011111111111111110000000000000000000111111111000000000000000000000000000000000000000000000001111111111111000000;
7'd51:player<=220'b0111111111111111100000001111100000000000000000000011111110000000111110000000001111110000111111111111111110000011111111111111111000000000000000001111111111100000000000000000000000000000000000000000000111111111111111100000;
7'd52:player<=220'b0111111111111111110000001111100000000000000000000111111110000000111111000000001111110000111111111111111110000011111111111111111100000000000000011111111111110000000000000000000000000000000000000000000111111111111111110000;
7'd53:player<=220'b0111111111111111110000001111100000000000000000000111111110000000011111000000001111100000111111111111111110000011111111111111111100000000000000011111111111111000000000000000000000000000000000000000001111111111111111111000;
7'd54:player<=220'b0111110000011111111000001111100000000000000000000111111110000000011111100000011111100000111111111111111100000011111111111111111110000000000000111111111111111000000000000000000000000000000000000000011111111000011111111000;
7'd55:player<=220'b0111110000000111111000001111100000000000000000001111111111000000011111100000011111000000111110000000000000000011111000000011111110000000000000111111000111111000000000000000000000000000000000000000011111100000000111111100;
7'd56:player<=220'b0111110000000111111000001111100000000000000000001111111111000000001111100000111111000000111110000000000000000011111000000001111110000000000000111110000011111100000000000000000000000000000000000000111111100000000011111100;
7'd57:player<=220'b0111110000000011111000001111100000000000000000001111101111000000001111110000111111000000111110000000000000000011111000000000111110000000000001111100000011111100000000000000000000000000000000000000111111000000000001111100;
7'd58:player<=220'b0111110000000011111000001111100000000000000000001111001111000000000111110000111110000000111110000000000000000011111000000000111110000000000001111100000001111100000000000000000000000000000000000000111110000000000001111110;
7'd59:player<=220'b0111110000000011111100001111100000000000000000011111001111100000000111111001111110000000111110000000000000000011111000000000111110000000000001111100000001111100000000000000000000000000000000000001111110000000000001111110;
7'd60:player<=220'b0111110000000011111000001111100000000000000000011111001111100000000011111001111100000000111110000000000000000011111000000001111110000000000000000000000001111100000000000000000000000000000000000001111110000000000000111110;
7'd61:player<=220'b0111110000000011111000001111100000000000000000011111000111100000000011111011111100000000111110000000000000000011111000000001111100000000000000000000000011111100000000000000000000000000000000000001111110000000000000111110;
7'd62:player<=220'b0111110000000111111000001111100000000000000000111110000111110000000011111111111000000000111111111111111100000011111000000011111100000000000000000000000011111000000000000000000000000000000000000001111110000000000000111110;
7'd63:player<=220'b0111110000001111111000001111100000000000000000111110000111110000000001111111111000000000111111111111111100000011111111111111111000000000000000000000000011111000000000000000000000000000000000000001111100000000000000111111;
7'd64:player<=220'b0111111111111111111000001111100000000000000000111110000111110000000001111111111000000000111111111111111100000011111111111111111000000000000000000000000111111000000000000000000000000000000000000001111100000000000000111111;
7'd65:player<=220'b0111111111111111110000001111100000000000000000111110000011110000000000111111110000000000111111111111111100000011111111111111100000000000000000000000001111110000000000000000000000000000000000000001111100000000000000111111;
7'd66:player<=220'b0111111111111111100000001111100000000000000001111100000011111000000000111111110000000000111111111111111100000011111111111111100000000000000000000000001111110000000000000000000000000000000000000001111100000000000000111111;
7'd67:player<=220'b0111111111111111100000001111100000000000000001111100000011111000000000111111100000000000111111111111111000000011111111111111110000000000000000000000011111100000000000001111111111111111100000000001111110000000000000111110;
7'd68:player<=220'b0111111111111110000000001111100000000000000001111100000011111000000000011111100000000000111110000000000000000011111111111111111000000000000000000000111111000000000000001111111111111111100000000001111110000000000000111110;
7'd69:player<=220'b0111111111111000000000001111100000000000000001111111111111111100000000011111100000000000111110000000000000000011111100000011111100000000000000000001111110000000000000001111111111111111100000000001111110000000000000111110;
7'd70:player<=220'b0111110000000000000000001111100000000000000011111111111111111100000000011111100000000000111110000000000000000011111000000001111100000000000000000011111100000000000000001111111111111111100000000001111110000000000001111110;
7'd71:player<=220'b0111110000000000000000001111100000000000000011111111111111111100000000011111100000000000111110000000000000000011111000000001111100000000000000000111111100000000000000001111111111111111100000000000111110000000000001111110;
7'd72:player<=220'b0111110000000000000000001111100000000000000011111111111111111100000000011111100000000000111110000000000000000011111000000001111110000000000000001111111000000000000000000000000000000000000000000000111111000000000001111110;
7'd73:player<=220'b0111110000000000000000001111100000000000000111111111111111111110000000011111100000000000111110000000000000000011111000000000111110000000000000001111110000000000000000000000000000000000000000000000111111000000000011111100;
7'd74:player<=220'b0111110000000000000000001111100000000000000111111000000001111110000000011111100000000000111110000000000000000011111000000000111110000000000000011111100000000000000000000000000000000000000000000000011111100000000111111100;
7'd75:player<=220'b0111110000000000000000001111111111111110000111110000000000111110000000011111100000000000111111000000000000000011111000000000111110000000000000111111000000000000000000000000000000000000000000000000011111110000001111111000;
7'd76:player<=220'b0111110000000000000000001111111111111111000111110000000000111111000000011111100000000000111111111111111110000011111000000000111111000000000001111111111111111100000000000000000000000000000000000000001111111111111111111000;
7'd77:player<=220'b0111110000000000000000001111111111111111001111110000000000111111000000011111100000000000111111111111111110000011111000000000111111000000000001111111111111111100000000000000000000000000000000000000001111111111111111110000;
7'd78:player<=220'b0111110000000000000000001111111111111111001111100000000000011111000000011111100000000000111111111111111110000011111000000000011111000000000001111111111111111100000000000000000000000000000000000000000111111111111111100000;
7'd79:player<=220'b0111110000000000000000001111111111111111001111100000000000011111000000011111100000000000111111111111111110000011111000000000011111000000000001111111111111111100000000000000000000000000000000000000000011111111111111000000;
7'd80:player<=220'b0111110000000000000000001111111111111111011111100000000000011111100000011111100000000000111111111111111110000011111000000000011111100000000001111111111111111100000000000000000000000000000000000000000000111111111110000000;
7'd81:player<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000;
        default:player<=0;
    endcase
end
endmodule

module WIN_LOGIC(clk_25M,win,win_adrs,win_sel);
input clk_25M;
input [1:0]win_sel;
output reg [0:219] win;
input [6:0] win_adrs;
always @(posedge clk_25M)
begin
    case(win_sel)
        2'b00:win<=0;
        2'b01:
        begin
            case(win_adrs)
                7'd00:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd01:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd02:win<=220'b0111111111111111100000000000000000000000000000011111111111111110000000000000000000000000000001111111111111111000000000011111111111111100000000000000000001111111111111111000000000000000000000000000000000011111111111111100;
                7'd03:win<=220'b0111111111111111110000000000000000000000000000011111111111111110000000000000000000000000000001111111111111111000000000011111111111111110000000000000000001111111111111111000000000000000000000000000000000011111111111111100;
                7'd04:win<=220'b0111111111111111110000000000000000000000000000111111111111111111000000000000000000000000000011111111111111110000000000011111111111111110000000000000000001111111111111111100000000000000000000000000000000011111111111111100;
                7'd05:win<=220'b0011111111111111110000000000000000000000000000111111111111111111000000000000000000000000000011111111111111110000000000011111111111111110000000000000000001111111111111111110000000000000000000000000000000011111111111111100;
                7'd06:win<=220'b0011111111111111110000000000000000000000000000111111111111111111000000000000000000000000000011111111111111110000000000011111111111111110000000000000000001111111111111111110000000000000000000000000000000011111111111111100;
                7'd07:win<=220'b0011111111111111111000000000000000000000000000111111111111111111000000000000000000000000000011111111111111110000000000011111111111111110000000000000000001111111111111111111000000000000000000000000000000011111111111111100;
                7'd08:win<=220'b0001111111111111111000000000000000000000000001111111111111111111100000000000000000000000000111111111111111100000000000011111111111111110000000000000000001111111111111111111100000000000000000000000000000011111111111111100;
                7'd09:win<=220'b0001111111111111111000000000000000000000000001111111111111111111100000000000000000000000000111111111111111100000000000011111111111111110000000000000000001111111111111111111100000000000000000000000000000011111111111111100;
                7'd10:win<=220'b0001111111111111111000000000000000000000000001111111111111111111100000000000000000000000000111111111111111100000000000011111111111111110000000000000000001111111111111111111110000000000000000000000000000011111111111111100;
                7'd11:win<=220'b0000111111111111111100000000000000000000000001111111111111111111110000000000000000000000001111111111111111000000000000011111111111111110000000000000000001111111111111111111111000000000000000000000000000011111111111111100;
                7'd12:win<=220'b0000111111111111111100000000000000000000000011111111111111111111110000000000000000000000001111111111111111000000000000011111111111111110000000000000000001111111111111111111111000000000000000000000000000011111111111111100;
                7'd13:win<=220'b0000111111111111111100000000000000000000000011111111111111111111110000000000000000000000001111111111111111000000000000011111111111111110000000000000000001111111111111111111111100000000000000000000000000011111111111111100;
                7'd14:win<=220'b0000111111111111111100000000000000000000000011111111111111111111110000000000000000000000001111111111111110000000000000011111111111111110000000000000000001111111111111111111111110000000000000000000000000011111111111111100;
                7'd15:win<=220'b0000011111111111111110000000000000000000000111111111111111111111111000000000000000000000011111111111111110000000000000011111111111111110000000000000000001111111111111111111111111000000000000000000000000011111111111111100;
                7'd16:win<=220'b0000011111111111111110000000000000000000000111111111111111111111111000000000000000000000011111111111111110000000000000011111111111111110000000000000000001111111111111111111111111000000000000000000000000011111111111111100;
                7'd17:win<=220'b0000011111111111111110000000000000000000000111111111111111111111111000000000000000000000011111111111111110000000000000011111111111111110000000000000000001111111111111111111111111100000000000000000000000011111111111111100;
                7'd18:win<=220'b0000001111111111111110000000000000000000000111111111111111111111111000000000000000000000011111111111111100000000000000011111111111111110000000000000000001111111111111111111111111110000000000000000000000011111111111111100;
                7'd19:win<=220'b0000001111111111111111000000000000000000001111111111111111111111111100000000000000000000111111111111111100000000000000011111111111111110000000000000000001111111111111111111111111110000000000000000000000011111111111111100;
                7'd20:win<=220'b0000001111111111111111000000000000000000001111111111111111111111111100000000000000000000111111111111111100000000000000011111111111111110000000000000000001111111111111111111111111111000000000000000000000011111111111111100;
                7'd21:win<=220'b0000000111111111111111000000000000000000001111111111111111111111111100000000000000000000111111111111111000000000000000011111111111111110000000000000000001111111111111111111111111111100000000000000000000011111111111111100;
                7'd22:win<=220'b0000000111111111111111000000000000000000001111111111111111111111111110000000000000000000111111111111111000000000000000011111111111111110000000000000000001111111111111111111111111111100000000000000000000011111111111111100;
                7'd23:win<=220'b0000000111111111111111100000000000000000011111111111110111111111111110000000000000000001111111111111111000000000000000011111111111111110000000000000000001111111111111111111111111111110000000000000000000011111111111111100;
                7'd24:win<=220'b0000000111111111111111100000000000000000011111111111110011111111111110000000000000000001111111111111110000000000000000011111111111111110000000000000000001111111111111111111111111111111000000000000000000011111111111111100;
                7'd25:win<=220'b0000000011111111111111100000000000000000011111111111110011111111111110000000000000000001111111111111110000000000000000011111111111111110000000000000000001111111111111111111111111111111000000000000000000011111111111111100;
                7'd26:win<=220'b0000000011111111111111110000000000000000011111111111110011111111111111000000000000000001111111111111110000000000000000011111111111111110000000000000000001111111111111111111111111111111100000000000000000011111111111111100;
                7'd27:win<=220'b0000000011111111111111110000000000000000111111111111100011111111111111000000000000000011111111111111110000000000000000011111111111111110000000000000000001111111111111111111111111111111110000000000000000011111111111111100;
                7'd28:win<=220'b0000000001111111111111110000000000000000111111111111100001111111111111000000000000000011111111111111100000000000000000011111111111111110000000000000000001111111111111110111111111111111110000000000000000011111111111111100;
                7'd29:win<=220'b0000000001111111111111110000000000000000111111111111100001111111111111000000000000000011111111111111100000000000000000011111111111111110000000000000000001111111111111110011111111111111111000000000000000011111111111111100;
                7'd30:win<=220'b0000000001111111111111111000000000000001111111111111100001111111111111100000000000000011111111111111100000000000000000011111111111111110000000000000000001111111111111110011111111111111111100000000000000011111111111111100;
                7'd31:win<=220'b0000000001111111111111111000000000000001111111111111000001111111111111100000000000000111111111111111000000000000000000011111111111111110000000000000000001111111111111110001111111111111111100000000000000011111111111111100;
                7'd32:win<=220'b0000000000111111111111111000000000000001111111111111000000111111111111100000000000000111111111111111000000000000000000011111111111111110000000000000000001111111111111110000111111111111111110000000000000011111111111111100;
                7'd33:win<=220'b0000000000111111111111111000000000000001111111111111000000111111111111100000000000000111111111111111000000000000000000011111111111111110000000000000000001111111111111110000111111111111111111000000000000011111111111111100;
                7'd34:win<=220'b0000000000111111111111111100000000000011111111111110000000111111111111110000000000000111111111111110000000000000000000011111111111111110000000000000000001111111111111110000011111111111111111100000000000011111111111111100;
                7'd35:win<=220'b0000000000011111111111111100000000000011111111111110000000011111111111110000000000001111111111111110000000000000000000011111111111111110000000000000000001111111111111110000001111111111111111100000000000011111111111111100;
                7'd36:win<=220'b0000000000011111111111111100000000000011111111111110000000011111111111110000000000001111111111111110000000000000000000011111111111111110000000000000000001111111111111110000001111111111111111110000000000011111111111111100;
                7'd37:win<=220'b0000000000011111111111111100000000000011111111111110000000011111111111111000000000001111111111111110000000000000000000011111111111111110000000000000000001111111111111110000000111111111111111111000000000011111111111111100;
                7'd38:win<=220'b0000000000001111111111111110000000000111111111111100000000011111111111111000000000001111111111111100000000000000000000011111111111111110000000000000000001111111111111110000000011111111111111111000000000011111111111111100;
                7'd39:win<=220'b0000000000001111111111111110000000000111111111111100000000001111111111111000000000011111111111111100000000000000000000011111111111111110000000000000000001111111111111110000000011111111111111111100000000011111111111111100;
                7'd40:win<=220'b0000000000001111111111111110000000000111111111111100000000001111111111111000000000011111111111111100000000000000000000011111111111111110000000000000000001111111111111110000000001111111111111111110000000011111111111111100;
                7'd41:win<=220'b0000000000001111111111111110000000000111111111111100000000001111111111111100000000011111111111111000000000000000000000011111111111111110000000000000000001111111111111110000000000111111111111111110000000011111111111111100;
                7'd42:win<=220'b0000000000000111111111111111000000001111111111111000000000001111111111111100000000011111111111111000000000000000000000011111111111111110000000000000000001111111111111110000000000111111111111111111000000011111111111111100;
                7'd43:win<=220'b0000000000000111111111111111000000001111111111111000000000000111111111111100000000111111111111111000000000000000000000011111111111111110000000000000000001111111111111110000000000011111111111111111100000011111111111111100;
                7'd44:win<=220'b0000000000000111111111111111000000001111111111111000000000000111111111111100000000111111111111110000000000000000000000011111111111111110000000000000000001111111111111110000000000001111111111111111100000011111111111111100;
                7'd45:win<=220'b0000000000000011111111111111000000011111111111111000000000000111111111111110000000111111111111110000000000000000000000011111111111111110000000000000000001111111111111110000000000001111111111111111110000011111111111111100;
                7'd46:win<=220'b0000000000000011111111111111100000011111111111110000000000000111111111111110000000111111111111110000000000000000000000011111111111111110000000000000000001111111111111110000000000000111111111111111111000011111111111111100;
                7'd47:win<=220'b0000000000000011111111111111100000011111111111110000000000000011111111111110000001111111111111110000000000000000000000011111111111111110000000000000000001111111111111110000000000000011111111111111111000011111111111111100;
                7'd48:win<=220'b0000000000000001111111111111100000011111111111110000000000000011111111111111000001111111111111100000000000000000000000011111111111111110000000000000000001111111111111110000000000000011111111111111111100011111111111111100;
                7'd49:win<=220'b0000000000000001111111111111100000111111111111110000000000000011111111111111000001111111111111100000000000000000000000011111111111111110000000000000000001111111111111110000000000000001111111111111111110011111111111111100;
                7'd50:win<=220'b0000000000000001111111111111110000111111111111100000000000000011111111111111000001111111111111100000000000000000000000011111111111111110000000000000000001111111111111110000000000000000111111111111111110011111111111111100;
                7'd51:win<=220'b0000000000000001111111111111110000111111111111100000000000000001111111111111000011111111111111000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000011111111111111111011111111111111100;
                7'd52:win<=220'b0000000000000000111111111111110000111111111111100000000000000001111111111111100011111111111111000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000011111111111111111111111111111111100;
                7'd53:win<=220'b0000000000000000111111111111110001111111111111100000000000000001111111111111100011111111111111000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000001111111111111111111111111111111100;
                7'd54:win<=220'b0000000000000000111111111111111001111111111111000000000000000000111111111111100011111111111110000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000111111111111111111111111111111100;
                7'd55:win<=220'b0000000000000000011111111111111001111111111111000000000000000000111111111111100111111111111110000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000111111111111111111111111111111100;
                7'd56:win<=220'b0000000000000000011111111111111001111111111111000000000000000000111111111111110111111111111110000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000011111111111111111111111111111100;
                7'd57:win<=220'b0000000000000000011111111111111011111111111110000000000000000000111111111111110111111111111110000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000001111111111111111111111111111100;
                7'd58:win<=220'b0000000000000000001111111111111111111111111110000000000000000000011111111111111111111111111100000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000001111111111111111111111111111100;
                7'd59:win<=220'b0000000000000000001111111111111111111111111110000000000000000000011111111111111111111111111100000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000111111111111111111111111111100;
                7'd60:win<=220'b0000000000000000001111111111111111111111111110000000000000000000011111111111111111111111111100000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000011111111111111111111111111100;
                7'd61:win<=220'b0000000000000000001111111111111111111111111100000000000000000000011111111111111111111111111000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000011111111111111111111111111100;
                7'd62:win<=220'b0000000000000000000111111111111111111111111100000000000000000000001111111111111111111111111000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000001111111111111111111111111100;
                7'd63:win<=220'b0000000000000000000111111111111111111111111100000000000000000000001111111111111111111111111000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000111111111111111111111111100;
                7'd64:win<=220'b0000000000000000000111111111111111111111111100000000000000000000001111111111111111111111110000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000111111111111111111111111100;
                7'd65:win<=220'b0000000000000000000011111111111111111111111000000000000000000000001111111111111111111111110000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000011111111111111111111111100;
                7'd66:win<=220'b0000000000000000000011111111111111111111111000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000001111111111111111111111100;
                7'd67:win<=220'b0000000000000000000011111111111111111111111000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000001111111111111111111111100;
                7'd68:win<=220'b0000000000000000000011111111111111111111111000000000000000000000000111111111111111111111100000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000111111111111111111111100;
                7'd69:win<=220'b0000000000000000000001111111111111111111110000000000000000000000000111111111111111111111100000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000011111111111111111111100;
                7'd70:win<=220'b0000000000000000000001111111111111111111110000000000000000000000000011111111111111111111100000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000011111111111111111111100;
                7'd71:win<=220'b0000000000000000000001111111111111111111110000000000000000000000000011111111111111111111000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000001111111111111111111100;
                7'd72:win<=220'b0000000000000000000000111111111111111111110000000000000000000000000011111111111111111111000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000111111111111111111100;
                7'd73:win<=220'b0000000000000000000000111111111111111111100000000000000000000000000001111111111111111111000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000011111111111111111100;
                7'd74:win<=220'b0000000000000000000000111111111111111111100000000000000000000000000001111111111111111111000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000011111111111111111100;
                7'd75:win<=220'b0000000000000000000000011111111111111111100000000000000000000000000001111111111111111110000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000001111111111111111100;
                7'd76:win<=220'b0000000000000000000000011111111111111111100000000000000000000000000001111111111111111110000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000000111111111111111100;
                7'd77:win<=220'b0000000000000000000000011111111111111111000000000000000000000000000000111111111111111110000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000000111111111111111100;
                7'd78:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd79:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd80:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd81:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd82:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd83:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd84:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd85:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd86:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd87:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd88:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd89:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd90:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd91:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd92:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd93:win<=220'b0000000000011111111111111111000000000000001111110000000000000000000000000000111111110000000001111111100000000000000111111100001111111111111111111111100000011111111111111111100000000000000000000000000000000000000000000000;
                7'd94:win<=220'b0000000000011111111111111111110000000000001111111000000000000000000000000000111111110000000001111111100000000000001111111100001111111111111111111111100000011111111111111111111100000000000000000000000000000011111110000000;
                7'd95:win<=220'b0000000000011111111111111111111100000000001111111000000000000000000000000000111111111000000000111111110000000000001111111000001111111111111111111111100000011111111111111111111110000000000000000000000000000011111110000000;
                7'd96:win<=220'b0000000000011111111111111111111110000000001111111000000000000000000000000001111111111000000000011111110000000000011111111000001111111111111111111111100000011111111111111111111111000000000000000000000000001111111110000000;
                7'd97:win<=220'b0000000000011111111111111111111111000000001111111000000000000000000000000001111111111000000000011111111000000000011111110000001111111111111111111111100000011111111111111111111111100000000000000000000000011111111110000000;
                7'd98:win<=220'b0000000000011111111111111111111111100000001111111000000000000000000000000001111111111100000000001111111000000000111111100000001111111111111111111111100000011111111111111111111111110000000000000000000001111111111110000000;
                7'd99:win<=220'b0000000000011111110000000011111111100000001111111000000000000000000000000011111111111100000000001111111100000000111111100000001111111000000000000000000000011111110000000001111111110000000000000000001111111111111110000000;
                7'd100:win<=220'b0000000000011111110000000000111111110000001111111000000000000000000000000011111111111100000000000111111100000001111111000000001111111000000000000000000000011111110000000000111111110000000000000000001111111111111110000000;
                7'd101:win<=220'b0000000000011111110000000000111111110000001111111000000000000000000000000111111101111110000000000111111110000001111111000000001111111000000000000000000000011111110000000000011111110000000000000000001111111111111110000000;
                7'd102:win<=220'b0000000000011111110000000000011111110000001111111000000000000000000000000111111001111110000000000011111110000011111110000000001111111000000000000000000000011111110000000000011111110000000000000000001111111011111110000000;
                7'd103:win<=220'b0000000000011111110000000000011111110000001111111000000000000000000000000111111001111110000000000011111111000011111110000000001111111000000000000000000000011111110000000000011111110000000000000000001111110011111110000000;
                7'd104:win<=220'b0000000000011111110000000000011111110000001111111000000000000000000000001111111000111111000000000001111111000111111100000000001111111000000000000000000000011111110000000000011111110000000000000000001111000011111110000000;
                7'd105:win<=220'b0000000000011111110000000000011111110000001111111000000000000000000000001111110000111111000000000001111111100111111100000000001111111000000000000000000000011111110000000000011111110000000000000000001000000011111110000000;
                7'd106:win<=220'b0000000000011111110000000000111111110000001111111000000000000000000000001111110000111111100000000000111111101111111000000000001111111100000000000000000000011111110000000000111111100000000000000000000000000011111110000000;
                7'd107:win<=220'b0000000000011111110000000001111111100000001111111000000000000000000000011111110000011111100000000000011111111111111000000000001111111111111111111110000000011111110000000011111111100000000000000000000000000011111110000000;
                7'd108:win<=220'b0000000000011111110000000011111111100000001111111000000000000000000000011111100000011111100000000000011111111111110000000000001111111111111111111110000000011111111111111111111111000000000000000000000000000011111110000000;
                7'd109:win<=220'b0000000000011111111111111111111111100000001111111000000000000000000000011111100000011111110000000000001111111111110000000000001111111111111111111110000000011111111111111111111100000000000000000000000000000011111110000000;
                7'd110:win<=220'b0000000000011111111111111111111111000000001111111000000000000000000000111111100000011111110000000000001111111111100000000000001111111111111111111110000000011111111111111111111000000000000000000000000000000011111110000000;
                7'd111:win<=220'b0000000000011111111111111111111110000000001111111000000000000000000000111111000000001111110000000000000111111111000000000000001111111111111111111110000000011111111111111111111100000000000000000000000000000011111110000000;
                7'd112:win<=220'b0000000000011111111111111111111100000000001111111000000000000000000001111111000000001111111000000000000111111111000000000000001111111100000000000000000000011111111111111111111110000000000000000000000000000011111110000000;
                7'd113:win<=220'b0000000000011111111111111111110000000000001111111000000000000000000001111111111111111111111000000000000011111110000000000000001111111000000000000000000000011111111111111111111111000000000000000000000000000011111110000000;
                7'd114:win<=220'b0000000000011111111111110000000000000000001111111000000000000000000001111111111111111111111000000000000011111110000000000000001111111000000000000000000000011111110000000001111111100000000000000000000000000011111110000000;
                7'd115:win<=220'b0000000000011111110000000000000000000000001111111000000000000000000011111111111111111111111100000000000011111110000000000000001111111000000000000000000000011111110000000000111111100000000000000000000000000011111110000000;
                7'd116:win<=220'b0000000000011111110000000000000000000000001111111000000000000000000011111111111111111111111100000000000011111110000000000000001111111000000000000000000000011111110000000000011111110000000000000000000000000011111110000000;
                7'd117:win<=220'b0000000000011111110000000000000000000000001111111000000000000000000011111111111111111111111110000000000011111110000000000000001111111000000000000000000000011111110000000000011111110000000000000000000000000011111110000000;
                7'd118:win<=220'b0000000000011111110000000000000000000000001111111000000000000000000111111111111111111111111110000000000011111110000000000000001111111000000000000000000000011111110000000000011111110000000000000000000000000011111110000000;
                7'd119:win<=220'b0000000000011111110000000000000000000000001111111000000000000000000111111100000000000011111110000000000011111110000000000000001111111000000000000000000000011111110000000000001111111000000000000000000000000011111110000000;
                7'd120:win<=220'b0000000000011111110000000000000000000000001111111111111111111100000111111100000000000001111111000000000011111110000000000000001111111100000000000000000000011111110000000000001111111000000000000000000000000011111110000000;
                7'd121:win<=220'b0000000000011111110000000000000000000000001111111111111111111110001111111000000000000001111111000000000011111110000000000000001111111111111111111111100000011111110000000000001111111000000000000000000000000011111110000000;
                7'd122:win<=220'b0000000000011111110000000000000000000000001111111111111111111110001111111000000000000001111111000000000011111110000000000000001111111111111111111111100000011111110000000000001111111000000000000000000000000011111110000000;
                7'd123:win<=220'b0000000000011111110000000000000000000000001111111111111111111110011111111000000000000000111111100000000011111110000000000000001111111111111111111111100000011111110000000000000111111100000000000000000000000011111110000000;
                7'd124:win<=220'b0000000000011111110000000000000000000000001111111111111111111110011111110000000000000000111111100000000011111110000000000000001111111111111111111111100000011111110000000000000111111100000000000000000000000011111110000000;
                7'd125:win<=220'b0000000000011111110000000000000000000000001111111111111111111110011111110000000000000000111111100000000011111110000000000000001111111111111111111111100000011111110000000000000111111100000000000000000000000011111110000000;
                7'd126:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd127:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            endcase
        end
        2'b10:
        begin
            case(win_adrs)
                7'd00:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd01:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd02:win<=220'b0111111111111111100000000000000000000000000000011111111111111110000000000000000000000000000001111111111111111000000000011111111111111100000000000000000001111111111111111000000000000000000000000000000000011111111111111100;
                7'd03:win<=220'b0111111111111111110000000000000000000000000000011111111111111110000000000000000000000000000001111111111111111000000000011111111111111110000000000000000001111111111111111000000000000000000000000000000000011111111111111100;
                7'd04:win<=220'b0111111111111111110000000000000000000000000000111111111111111111000000000000000000000000000011111111111111110000000000011111111111111110000000000000000001111111111111111100000000000000000000000000000000011111111111111100;
                7'd05:win<=220'b0011111111111111110000000000000000000000000000111111111111111111000000000000000000000000000011111111111111110000000000011111111111111110000000000000000001111111111111111110000000000000000000000000000000011111111111111100;
                7'd06:win<=220'b0011111111111111110000000000000000000000000000111111111111111111000000000000000000000000000011111111111111110000000000011111111111111110000000000000000001111111111111111110000000000000000000000000000000011111111111111100;
                7'd07:win<=220'b0011111111111111111000000000000000000000000000111111111111111111000000000000000000000000000011111111111111110000000000011111111111111110000000000000000001111111111111111111000000000000000000000000000000011111111111111100;
                7'd08:win<=220'b0001111111111111111000000000000000000000000001111111111111111111100000000000000000000000000111111111111111100000000000011111111111111110000000000000000001111111111111111111100000000000000000000000000000011111111111111100;
                7'd09:win<=220'b0001111111111111111000000000000000000000000001111111111111111111100000000000000000000000000111111111111111100000000000011111111111111110000000000000000001111111111111111111100000000000000000000000000000011111111111111100;
                7'd10:win<=220'b0001111111111111111000000000000000000000000001111111111111111111100000000000000000000000000111111111111111100000000000011111111111111110000000000000000001111111111111111111110000000000000000000000000000011111111111111100;
                7'd11:win<=220'b0000111111111111111100000000000000000000000001111111111111111111110000000000000000000000001111111111111111000000000000011111111111111110000000000000000001111111111111111111111000000000000000000000000000011111111111111100;
                7'd12:win<=220'b0000111111111111111100000000000000000000000011111111111111111111110000000000000000000000001111111111111111000000000000011111111111111110000000000000000001111111111111111111111000000000000000000000000000011111111111111100;
                7'd13:win<=220'b0000111111111111111100000000000000000000000011111111111111111111110000000000000000000000001111111111111111000000000000011111111111111110000000000000000001111111111111111111111100000000000000000000000000011111111111111100;
                7'd14:win<=220'b0000111111111111111100000000000000000000000011111111111111111111110000000000000000000000001111111111111110000000000000011111111111111110000000000000000001111111111111111111111110000000000000000000000000011111111111111100;
                7'd15:win<=220'b0000011111111111111110000000000000000000000111111111111111111111111000000000000000000000011111111111111110000000000000011111111111111110000000000000000001111111111111111111111111000000000000000000000000011111111111111100;
                7'd16:win<=220'b0000011111111111111110000000000000000000000111111111111111111111111000000000000000000000011111111111111110000000000000011111111111111110000000000000000001111111111111111111111111000000000000000000000000011111111111111100;
                7'd17:win<=220'b0000011111111111111110000000000000000000000111111111111111111111111000000000000000000000011111111111111110000000000000011111111111111110000000000000000001111111111111111111111111100000000000000000000000011111111111111100;
                7'd18:win<=220'b0000001111111111111110000000000000000000000111111111111111111111111000000000000000000000011111111111111100000000000000011111111111111110000000000000000001111111111111111111111111110000000000000000000000011111111111111100;
                7'd19:win<=220'b0000001111111111111111000000000000000000001111111111111111111111111100000000000000000000111111111111111100000000000000011111111111111110000000000000000001111111111111111111111111110000000000000000000000011111111111111100;
                7'd20:win<=220'b0000001111111111111111000000000000000000001111111111111111111111111100000000000000000000111111111111111100000000000000011111111111111110000000000000000001111111111111111111111111111000000000000000000000011111111111111100;
                7'd21:win<=220'b0000000111111111111111000000000000000000001111111111111111111111111100000000000000000000111111111111111000000000000000011111111111111110000000000000000001111111111111111111111111111100000000000000000000011111111111111100;
                7'd22:win<=220'b0000000111111111111111000000000000000000001111111111111111111111111110000000000000000000111111111111111000000000000000011111111111111110000000000000000001111111111111111111111111111100000000000000000000011111111111111100;
                7'd23:win<=220'b0000000111111111111111100000000000000000011111111111110111111111111110000000000000000001111111111111111000000000000000011111111111111110000000000000000001111111111111111111111111111110000000000000000000011111111111111100;
                7'd24:win<=220'b0000000111111111111111100000000000000000011111111111110011111111111110000000000000000001111111111111110000000000000000011111111111111110000000000000000001111111111111111111111111111111000000000000000000011111111111111100;
                7'd25:win<=220'b0000000011111111111111100000000000000000011111111111110011111111111110000000000000000001111111111111110000000000000000011111111111111110000000000000000001111111111111111111111111111111000000000000000000011111111111111100;
                7'd26:win<=220'b0000000011111111111111110000000000000000011111111111110011111111111111000000000000000001111111111111110000000000000000011111111111111110000000000000000001111111111111111111111111111111100000000000000000011111111111111100;
                7'd27:win<=220'b0000000011111111111111110000000000000000111111111111100011111111111111000000000000000011111111111111110000000000000000011111111111111110000000000000000001111111111111111111111111111111110000000000000000011111111111111100;
                7'd28:win<=220'b0000000001111111111111110000000000000000111111111111100001111111111111000000000000000011111111111111100000000000000000011111111111111110000000000000000001111111111111110111111111111111110000000000000000011111111111111100;
                7'd29:win<=220'b0000000001111111111111110000000000000000111111111111100001111111111111000000000000000011111111111111100000000000000000011111111111111110000000000000000001111111111111110011111111111111111000000000000000011111111111111100;
                7'd30:win<=220'b0000000001111111111111111000000000000001111111111111100001111111111111100000000000000011111111111111100000000000000000011111111111111110000000000000000001111111111111110011111111111111111100000000000000011111111111111100;
                7'd31:win<=220'b0000000001111111111111111000000000000001111111111111000001111111111111100000000000000111111111111111000000000000000000011111111111111110000000000000000001111111111111110001111111111111111100000000000000011111111111111100;
                7'd32:win<=220'b0000000000111111111111111000000000000001111111111111000000111111111111100000000000000111111111111111000000000000000000011111111111111110000000000000000001111111111111110000111111111111111110000000000000011111111111111100;
                7'd33:win<=220'b0000000000111111111111111000000000000001111111111111000000111111111111100000000000000111111111111111000000000000000000011111111111111110000000000000000001111111111111110000111111111111111111000000000000011111111111111100;
                7'd34:win<=220'b0000000000111111111111111100000000000011111111111110000000111111111111110000000000000111111111111110000000000000000000011111111111111110000000000000000001111111111111110000011111111111111111100000000000011111111111111100;
                7'd35:win<=220'b0000000000011111111111111100000000000011111111111110000000011111111111110000000000001111111111111110000000000000000000011111111111111110000000000000000001111111111111110000001111111111111111100000000000011111111111111100;
                7'd36:win<=220'b0000000000011111111111111100000000000011111111111110000000011111111111110000000000001111111111111110000000000000000000011111111111111110000000000000000001111111111111110000001111111111111111110000000000011111111111111100;
                7'd37:win<=220'b0000000000011111111111111100000000000011111111111110000000011111111111111000000000001111111111111110000000000000000000011111111111111110000000000000000001111111111111110000000111111111111111111000000000011111111111111100;
                7'd38:win<=220'b0000000000001111111111111110000000000111111111111100000000011111111111111000000000001111111111111100000000000000000000011111111111111110000000000000000001111111111111110000000011111111111111111000000000011111111111111100;
                7'd39:win<=220'b0000000000001111111111111110000000000111111111111100000000001111111111111000000000011111111111111100000000000000000000011111111111111110000000000000000001111111111111110000000011111111111111111100000000011111111111111100;
                7'd40:win<=220'b0000000000001111111111111110000000000111111111111100000000001111111111111000000000011111111111111100000000000000000000011111111111111110000000000000000001111111111111110000000001111111111111111110000000011111111111111100;
                7'd41:win<=220'b0000000000001111111111111110000000000111111111111100000000001111111111111100000000011111111111111000000000000000000000011111111111111110000000000000000001111111111111110000000000111111111111111110000000011111111111111100;
                7'd42:win<=220'b0000000000000111111111111111000000001111111111111000000000001111111111111100000000011111111111111000000000000000000000011111111111111110000000000000000001111111111111110000000000111111111111111111000000011111111111111100;
                7'd43:win<=220'b0000000000000111111111111111000000001111111111111000000000000111111111111100000000111111111111111000000000000000000000011111111111111110000000000000000001111111111111110000000000011111111111111111100000011111111111111100;
                7'd44:win<=220'b0000000000000111111111111111000000001111111111111000000000000111111111111100000000111111111111110000000000000000000000011111111111111110000000000000000001111111111111110000000000001111111111111111100000011111111111111100;
                7'd45:win<=220'b0000000000000011111111111111000000011111111111111000000000000111111111111110000000111111111111110000000000000000000000011111111111111110000000000000000001111111111111110000000000001111111111111111110000011111111111111100;
                7'd46:win<=220'b0000000000000011111111111111100000011111111111110000000000000111111111111110000000111111111111110000000000000000000000011111111111111110000000000000000001111111111111110000000000000111111111111111111000011111111111111100;
                7'd47:win<=220'b0000000000000011111111111111100000011111111111110000000000000011111111111110000001111111111111110000000000000000000000011111111111111110000000000000000001111111111111110000000000000011111111111111111000011111111111111100;
                7'd48:win<=220'b0000000000000001111111111111100000011111111111110000000000000011111111111111000001111111111111100000000000000000000000011111111111111110000000000000000001111111111111110000000000000011111111111111111100011111111111111100;
                7'd49:win<=220'b0000000000000001111111111111100000111111111111110000000000000011111111111111000001111111111111100000000000000000000000011111111111111110000000000000000001111111111111110000000000000001111111111111111110011111111111111100;
                7'd50:win<=220'b0000000000000001111111111111110000111111111111100000000000000011111111111111000001111111111111100000000000000000000000011111111111111110000000000000000001111111111111110000000000000000111111111111111110011111111111111100;
                7'd51:win<=220'b0000000000000001111111111111110000111111111111100000000000000001111111111111000011111111111111000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000011111111111111111011111111111111100;
                7'd52:win<=220'b0000000000000000111111111111110000111111111111100000000000000001111111111111100011111111111111000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000011111111111111111111111111111111100;
                7'd53:win<=220'b0000000000000000111111111111110001111111111111100000000000000001111111111111100011111111111111000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000001111111111111111111111111111111100;
                7'd54:win<=220'b0000000000000000111111111111111001111111111111000000000000000000111111111111100011111111111110000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000111111111111111111111111111111100;
                7'd55:win<=220'b0000000000000000011111111111111001111111111111000000000000000000111111111111100111111111111110000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000111111111111111111111111111111100;
                7'd56:win<=220'b0000000000000000011111111111111001111111111111000000000000000000111111111111110111111111111110000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000011111111111111111111111111111100;
                7'd57:win<=220'b0000000000000000011111111111111011111111111110000000000000000000111111111111110111111111111110000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000001111111111111111111111111111100;
                7'd58:win<=220'b0000000000000000001111111111111111111111111110000000000000000000011111111111111111111111111100000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000001111111111111111111111111111100;
                7'd59:win<=220'b0000000000000000001111111111111111111111111110000000000000000000011111111111111111111111111100000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000111111111111111111111111111100;
                7'd60:win<=220'b0000000000000000001111111111111111111111111110000000000000000000011111111111111111111111111100000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000011111111111111111111111111100;
                7'd61:win<=220'b0000000000000000001111111111111111111111111100000000000000000000011111111111111111111111111000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000011111111111111111111111111100;
                7'd62:win<=220'b0000000000000000000111111111111111111111111100000000000000000000001111111111111111111111111000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000001111111111111111111111111100;
                7'd63:win<=220'b0000000000000000000111111111111111111111111100000000000000000000001111111111111111111111111000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000111111111111111111111111100;
                7'd64:win<=220'b0000000000000000000111111111111111111111111100000000000000000000001111111111111111111111110000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000111111111111111111111111100;
                7'd65:win<=220'b0000000000000000000011111111111111111111111000000000000000000000001111111111111111111111110000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000011111111111111111111111100;
                7'd66:win<=220'b0000000000000000000011111111111111111111111000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000001111111111111111111111100;
                7'd67:win<=220'b0000000000000000000011111111111111111111111000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000001111111111111111111111100;
                7'd68:win<=220'b0000000000000000000011111111111111111111111000000000000000000000000111111111111111111111100000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000111111111111111111111100;
                7'd69:win<=220'b0000000000000000000001111111111111111111110000000000000000000000000111111111111111111111100000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000011111111111111111111100;
                7'd70:win<=220'b0000000000000000000001111111111111111111110000000000000000000000000011111111111111111111100000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000011111111111111111111100;
                7'd71:win<=220'b0000000000000000000001111111111111111111110000000000000000000000000011111111111111111111000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000001111111111111111111100;
                7'd72:win<=220'b0000000000000000000000111111111111111111110000000000000000000000000011111111111111111111000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000111111111111111111100;
                7'd73:win<=220'b0000000000000000000000111111111111111111100000000000000000000000000001111111111111111111000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000011111111111111111100;
                7'd74:win<=220'b0000000000000000000000111111111111111111100000000000000000000000000001111111111111111111000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000011111111111111111100;
                7'd75:win<=220'b0000000000000000000000011111111111111111100000000000000000000000000001111111111111111110000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000001111111111111111100;
                7'd76:win<=220'b0000000000000000000000011111111111111111100000000000000000000000000001111111111111111110000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000000111111111111111100;
                7'd77:win<=220'b0000000000000000000000011111111111111111000000000000000000000000000000111111111111111110000000000000000000000000000000011111111111111110000000000000000001111111111111110000000000000000000000000000000000111111111111111100;
                7'd78:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd79:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd80:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd81:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd82:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd83:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd84:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd85:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd86:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd87:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd88:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd89:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd90:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd91:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd92:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd93:win<=220'b0000000000011111111111111111000000000000001111110000000000000000000000000000111111110000000001111111100000000000000111111100001111111111111111111111100000011111111111111111100000000000000000000000000000000000000000000000;
                7'd94:win<=220'b0000000000011111111111111111110000000000001111111000000000000000000000000000111111110000000001111111100000000000001111111100001111111111111111111111100000011111111111111111111100000000000000000000000111111110000000000000;
                7'd95:win<=220'b0000000000011111111111111111111100000000001111111000000000000000000000000000111111111000000000111111110000000000001111111000001111111111111111111111100000011111111111111111111110000000000000000000111111111111110000000000;
                7'd96:win<=220'b0000000000011111111111111111111110000000001111111000000000000000000000000001111111111000000000011111110000000000011111111000001111111111111111111111100000011111111111111111111111000000000000000011111111111111111100000000;
                7'd97:win<=220'b0000000000011111111111111111111111000000001111111000000000000000000000000001111111111000000000011111111000000000011111110000001111111111111111111111100000011111111111111111111111100000000000000111111111111111111110000000;
                7'd98:win<=220'b0000000000011111111111111111111111100000001111111000000000000000000000000001111111111100000000001111111000000000111111100000001111111111111111111111100000011111111111111111111111110000000000001111111111111111111111000000;
                7'd99:win<=220'b0000000000011111110000000011111111100000001111111000000000000000000000000011111111111100000000001111111100000000111111100000001111111000000000000000000000011111110000000001111111110000000000001111111111111111111111000000;
                7'd100:win<=220'b0000000000011111110000000000111111110000001111111000000000000000000000000011111111111100000000000111111100000001111111000000001111111000000000000000000000011111110000000000111111110000000000111111111000000111111111000000;
                7'd101:win<=220'b0000000000011111110000000000111111110000001111111000000000000000000000000111111101111110000000000111111110000001111111000000001111111000000000000000000000011111110000000000011111110000000000111111110000000011111111000000;
                7'd102:win<=220'b0000000000011111110000000000011111110000001111111000000000000000000000000111111001111110000000000011111110000011111110000000001111111000000000000000000000011111110000000000011111110000000000111111100000000011111111000000;
                7'd103:win<=220'b0000000000011111110000000000011111110000001111111000000000000000000000000111111001111110000000000011111111000011111110000000001111111000000000000000000000011111110000000000011111110000000001111111100000000001111111000000;
                7'd104:win<=220'b0000000000011111110000000000011111110000001111111000000000000000000000001111111000111111000000000001111111000111111100000000001111111000000000000000000000011111110000000000011111110000000001111111000000000001111111000000;
                7'd105:win<=220'b0000000000011111110000000000011111110000001111111000000000000000000000001111110000111111000000000001111111100111111100000000001111111000000000000000000000011111110000000000011111110000000000000000000000000011111111000000;
                7'd106:win<=220'b0000000000011111110000000000111111110000001111111000000000000000000000001111110000111111100000000000111111101111111000000000001111111100000000000000000000011111110000000000111111100000000000000000000000000011111111000000;
                7'd107:win<=220'b0000000000011111110000000001111111100000001111111000000000000000000000011111110000011111100000000000011111111111111000000000001111111111111111111110000000011111110000000011111111100000000000000000000000000111111110000000;
                7'd108:win<=220'b0000000000011111110000000011111111100000001111111000000000000000000000011111100000011111100000000000011111111111110000000000001111111111111111111110000000011111111111111111111111000000000000000000000000000111111110000000;
                7'd109:win<=220'b0000000000011111111111111111111111100000001111111000000000000000000000011111100000011111110000000000001111111111110000000000001111111111111111111110000000011111111111111111111100000000000000000000000000001111111100000000;
                7'd110:win<=220'b0000000000011111111111111111111111000000001111111000000000000000000000111111100000011111110000000000001111111111100000000000001111111111111111111110000000011111111111111111111000000000000000000000000000111111111000000000;
                7'd111:win<=220'b0000000000011111111111111111111110000000001111111000000000000000000000111111000000001111110000000000000111111111000000000000001111111111111111111110000000011111111111111111111100000000000000000000000001111111110000000000;
                7'd112:win<=220'b0000000000011111111111111111111100000000001111111000000000000000000001111111000000001111111000000000000111111111000000000000001111111100000000000000000000011111111111111111111110000000000000000000000011111111100000000000;
                7'd113:win<=220'b0000000000011111111111111111110000000000001111111000000000000000000001111111111111111111111000000000000011111110000000000000001111111000000000000000000000011111111111111111111111000000000000000000001111111111000000000000;
                7'd114:win<=220'b0000000000011111111111110000000000000000001111111000000000000000000001111111111111111111111000000000000011111110000000000000001111111000000000000000000000011111110000000001111111100000000000000000011111111110000000000000;
                7'd115:win<=220'b0000000000011111110000000000000000000000001111111000000000000000000011111111111111111111111100000000000011111110000000000000001111111000000000000000000000011111110000000000111111100000000000000000111111111000000000000000;
                7'd116:win<=220'b0000000000011111110000000000000000000000001111111000000000000000000011111111111111111111111100000000000011111110000000000000001111111000000000000000000000011111110000000000011111110000000000000001111111110000000000000000;
                7'd117:win<=220'b0000000000011111110000000000000000000000001111111000000000000000000011111111111111111111111110000000000011111110000000000000001111111000000000000000000000011111110000000000011111110000000000000111111111100000000000000000;
                7'd118:win<=220'b0000000000011111110000000000000000000000001111111000000000000000000111111111111111111111111110000000000011111110000000000000001111111000000000000000000000011111110000000000011111110000000000001111111110000000000000000000;
                7'd119:win<=220'b0000000000011111110000000000000000000000001111111000000000000000000111111100000000000011111110000000000011111110000000000000001111111000000000000000000000011111110000000000001111111000000000011111111100000000000000000000;
                7'd120:win<=220'b0000000000011111110000000000000000000000001111111111111111111100000111111100000000000001111111000000000011111110000000000000001111111100000000000000000000011111110000000000001111111000000001111111111111111111111111100000;
                7'd121:win<=220'b0000000000011111110000000000000000000000001111111111111111111110001111111000000000000001111111000000000011111110000000000000001111111111111111111111100000011111110000000000001111111000000001111111111111111111111111100000;
                7'd122:win<=220'b0000000000011111110000000000000000000000001111111111111111111110001111111000000000000001111111000000000011111110000000000000001111111111111111111111100000011111110000000000001111111000000011111111111111111111111111100000;
                7'd123:win<=220'b0000000000011111110000000000000000000000001111111111111111111110011111111000000000000000111111100000000011111110000000000000001111111111111111111111100000011111110000000000000111111100000011111111111111111111111111100000;
                7'd124:win<=220'b0000000000011111110000000000000000000000001111111111111111111110011111110000000000000000111111100000000011111110000000000000001111111111111111111111100000011111110000000000000111111100000011111111111111111111111111100000;
                7'd125:win<=220'b0000000000011111110000000000000000000000001111111111111111111110011111110000000000000000111111100000000011111110000000000000001111111111111111111111100000011111110000000000000111111100000000000000000000000000000000000000;
                7'd126:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                7'd127:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            endcase
        end
        2'b11:
        begin
            case(win_adrs)
            7'd00:win <=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            7'd01:win <=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            7'd02:win <=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            7'd03:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd04:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd05:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd06:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd07:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd08:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd09:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd10:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd11:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd12:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd13:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd14:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd15:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd16:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd17:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd18:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd19:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd20:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd21:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd22:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd23:win <=220'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000;
            7'd24:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd25:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd26:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd27:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd28:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd29:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd30:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd31:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd32:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd33:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd34:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd35:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd36:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd37:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd38:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd39:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd40:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd41:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd42:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd43:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd44:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd45:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd46:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd47:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd48:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd49:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd50:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd51:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000;
            7'd52:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd53:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd54:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd55:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd56:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd57:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd58:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd59:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd60:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd61:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd62:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd63:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd64:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd65:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd66:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd67:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd68:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd69:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd70:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd71:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000;
            7'd72:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd73:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd74:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd75:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd76:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd77:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd78:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd79:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd80:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd81:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd82:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd83:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd84:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd85:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd86:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd87:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd88:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd89:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd90:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd91:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd92:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd93:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd94:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd95:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd96:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd97:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd98:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd99:win <=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd100:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd101:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            7'd102:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000;
            7'd103:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd104:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd105:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd106:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd107:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd108:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd109:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd110:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd111:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd112:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd113:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd114:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd115:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd116:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd117:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd118:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd119:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd120:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd121:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd122:win<=220'b0000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000;
            7'd123:win<=220'b0000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111110000;
            7'd124:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            7'd125:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            7'd126:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            7'd127:win<=220'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            endcase
        end
    endcase
end
endmodule
// Clock Division for 100MHz
module CLK_10Hz(clk_in,clk_out);
input clk_in;
output reg clk_out=0;
integer i;
always @(posedge clk_in)
begin
    if(i==4999999)
    begin
        clk_out<=~clk_out;
        i<=0;
    end
    else
        i<=i+1;
end
endmodule
