// Adding Reset logic to score 
module DINO_GAME(sys_clk,clk_25M,clk_100,hcount,vcount,jump,red,green,blue,rst_dino);
input sys_clk,rst_dino;
input jump;
output [3:0] red,green,blue;
input [9:0] hcount,vcount;
input clk_25M,clk_100;
wire [63:0] dino_data;
wire [79:0] obstacle_data;
wire [0:399] title;
wire [0:99] score_t;
wire [5:0] title_adrs;
wire [6:0] obstacle_adrs;
wire [9:0] dino_pos=200;
wire [5:0] dino_adrs;
wire [9:0] v_dino_pos;
wire [9:0] obstacle_pos;
wire [9:0] v_obstacle_pos=435;
wire [5:0] go_adrs;
wire [0:235] game_over;
wire reset,set1;
//// Stop Logic
reg stop=0;
wire [4:0] score_adrs;
wire [0:19] score1,score2,score3,score4;
always @(posedge clk_25M)
begin
    if((obstacle_pos>=dino_pos-50 && obstacle_pos<=dino_pos+45 && v_dino_pos>=485 && v_dino_pos<=515 )||(obstacle_pos>=dino_pos+10 && obstacle_pos<=dino_pos+40 && v_dino_pos>=440 && v_dino_pos<=515))// 70 is width of the Obstacle
    begin
        stop<=1;
    end
    else
        stop<=0;
end
assign stop_temp=stop;
assign reset=(set1&jump)|rst_dino;

wire [3:0] bcd3,bcd2,bcd1,bcd0;
wire [15:0] bcd;
SCORE Score_counter(sys_clk,bcd,stop_temp,reset);
assign bcd3=bcd[15:12];
assign bcd2=bcd[11:8];
assign bcd1=bcd[7:4];
assign bcd0=bcd[3:0];
DINO_DATA Data(clk_25M,dino_data,dino_adrs,title_adrs,obstacle_data,obstacle_adrs,title,score_adrs,score_t,go_adrs,game_over);
DISP_WRITE_DINO Writing(clk_25M,hcount,vcount,dino_pos,v_dino_pos,obstacle_pos,v_obstacle_pos,dino_data,dino_adrs,obstacle_data,obstacle_adrs,title,title_adrs,score1,score2,score3,score4,score_t,score_adrs,stop_temp,go_adrs,game_over,red,green,blue);
JUMP_DINO Jump(clk_100,reset,jump,stop_temp,v_dino_pos);
MOVE_OBSTACLE Move(clk_100,reset,jump,stop_temp,obstacle_pos,set1);
SCORE_DATA Score1(clk_25M,bcd0,score1,score_adrs);
SCORE_DATA Score2(clk_25M,bcd1,score2,score_adrs);
SCORE_DATA Score3(clk_25M,bcd2,score3,score_adrs);
SCORE_DATA Score4(clk_25M,bcd3,score4,score_adrs);
endmodule
module DISP_WRITE_DINO(clk_25M,hcount,vcount,dino_pos,v_dino_pos,obstacle_pos,v_obstacle_pos,dino_data,dino_adrs,obstacle_data,obstacle_adrs,title,title_adrs,score1,score2,score3,score4,score_t,score_adrs,stop_temp,go_adrs,game_over,red,green,blue);
input clk_25M,stop_temp;
input [9:0] hcount,vcount,v_dino_pos,dino_pos,obstacle_pos,v_obstacle_pos;
input [63:0] dino_data;
input [79:0] obstacle_data;
input [0:399] title;
input [0:19] score1;
input [0:19] score2;
input [0:19] score3;
input [0:19] score4;
input [0:99] score_t;
input [0:235] game_over;
output reg [4:0] score_adrs;
output reg [6:0] obstacle_adrs;
output reg [5:0] dino_adrs,go_adrs;
output reg [5:0] title_adrs;
output reg [3:0] red,green,blue;
always @(posedge clk_25M)
begin
    if((hcount>=144 && hcount<=784) && (vcount>=35 && vcount<=521))
        begin
            obstacle_adrs<=vcount-v_obstacle_pos;
            dino_adrs<=vcount-v_dino_pos;
            title_adrs<=vcount-50;
            score_adrs<=vcount-110;
            go_adrs<=vcount-263;
            if((hcount>=dino_pos && hcount<=dino_pos+64) && (vcount>=v_dino_pos-64 && vcount<=v_dino_pos)&&(dino_data[hcount-dino_pos]==1))
            begin
                {red,green,blue}<={4'b1111,4'b1111,4'b1111};
            end
            else if((hcount>=obstacle_pos && hcount<=obstacle_pos+60) && (vcount>=v_obstacle_pos && vcount<=v_obstacle_pos+80)&&(obstacle_data[hcount-obstacle_pos]==1))
            begin
                {red,green,blue}<={4'b0001,4'b1001,4'b0100};
            end
            else if((hcount>=264 && hcount<=664) && (vcount>=50 && vcount<=100)&&(title[hcount-264]==1))
            begin
                {red,green,blue}<={4'b0001,4'b1001,4'b1011};
            end
            else if((hcount>=750 && hcount<=770) && (vcount>=110 && vcount<=142)&&(score1[hcount-750]==1))
            begin
                {red,green,blue}<={4'b1011,4'b1011,4'b0100};
            end
            else if((hcount>=730 && hcount<=750) && (vcount>=110 && vcount<=142)&&(score2[hcount-730]==1))
            begin
                {red,green,blue}<={4'b1011,4'b1011,4'b0100};
            end
            else if((hcount>=710 && hcount<=730) && (vcount>=110 && vcount<=142)&&(score3[hcount-710]==1))
            begin
                {red,green,blue}<={4'b1011,4'b1011,4'b0100};
            end
            else if((hcount>=690 && hcount<=710) && (vcount>=110 && vcount<=142)&&(score4[hcount-690]==1))
            begin
                {red,green,blue}<={4'b1011,4'b1011,4'b0100};
            end
            else if((hcount>=590 && hcount<=689) && (vcount>=110 && vcount<=142)&&(score_t[hcount-590]==1))
            begin
                {red,green,blue}<={4'b1011,4'b1011,4'b0100};
            end
            else if((hcount>=346 && hcount<=582) && (vcount>=263 && vcount<=327)&&(game_over[hcount-346]==1)&& stop_temp)
            begin
                {red,green,blue}<={4'b1110,4'b0001,4'b0001};
            end
            else
                {red,green,blue}<={4'b0000,4'b0000,4'b0000}; 
        end
    else
        begin
            {red,green,blue}<={4'b0000,4'b0000,4'b0000};   
        end
end
endmodule

// Obstacle Moving Logic
module MOVE_OBSTACLE(clk_100,reset,jump,stop_temp,obstacle_pos,set1);
input clk_100,reset,jump,stop_temp;
output reg [9:0] obstacle_pos=600;
output reg  set1;
always @(posedge clk_100)
begin
    if(reset)
    begin
        obstacle_pos<=744;
        set1<=1;
    end
    else
    begin
        if(stop_temp)
        begin
            if(jump)
            begin
                set1<=1;
                obstacle_pos<=obstacle_pos;
                //block2<=block2;
            end
            else
            begin
                set1<=0;
                obstacle_pos<=obstacle_pos;
            end
        end
        else
        begin
            set1<=0;
            if(obstacle_pos==104)
                obstacle_pos<=784;
            else
                obstacle_pos<=obstacle_pos-1;
        end
    end
end
endmodule

// Dino Jumping Logic
module JUMP_DINO(clk_100,reset,jump,stop_temp,v_dino_pos);
input clk_100,jump,reset,stop_temp;
output reg [9:0]v_dino_pos=515;
reg temp=0;
always @(posedge clk_100)
begin
        if(reset)
            temp<=0;
        else if(v_dino_pos==350)
            temp<=0;
        else if(jump)
            if(v_dino_pos==515)
                temp<=jump;
            else
                temp<=temp;
        else
            temp<=temp;
end
always @(posedge clk_100)
begin
    if(reset)
        v_dino_pos<=515;
	else if(stop_temp)
        v_dino_pos<=v_dino_pos;
	else
	begin
		if(temp)
		begin
		  if(v_dino_pos>300)
			v_dino_pos<=v_dino_pos-1;
	      else
	        v_dino_pos<=v_dino_pos;
	    end
		else
	    begin
			if(v_dino_pos<515)
				v_dino_pos<=v_dino_pos+1;
			else
				v_dino_pos<=v_dino_pos;
	    end
	end
end
endmodule

module SCORE(clk,score,stop_temp,reset);
input clk,reset,stop_temp;
output [15:0] score;
reg clk_div;
integer i;
integer div;
reg [13:0] bin=0;
always @(posedge clk)
begin
    if(i==div)
    begin
        clk_div<=~clk_div;
        i<=0;
    end
    else
        i<=i+1;
end
always @(posedge clk)
begin
    if(bin <15)
        div<=49999999;
    else if( bin>=15 && bin <=30)
        div<=25999999;
    else if( bin>30 && bin <=50)
        div<=12599999;
    else if( bin>50 && bin <=100)
        div<=10000000;
    else if( bin>100 && bin <=1000)
        div<=4999999;
    else if( bin>1000 && bin <10000)
        div<=2599999;
    else
        div<=div;
end
always @(posedge clk_div, posedge reset)
begin
    if(reset)
        bin<=0;
    else if(stop_temp)
        bin<=bin;
    else
        bin<=bin+1;
end
BIN_BCD Binary_BCD(clk,bin,score);
endmodule
module BIN_BCD(
input clk,
input [13:0]bin,
output reg [15:0]bcd
);
reg [3:0]count=0;
reg [15:0] bcd_temp=0;
reg reset=0;
always@(posedge clk)
if(reset) begin
    bcd_temp=0;
    count=0;
    reset=0;
end
else if(count<=13)
begin
    if(bcd_temp[3:0]>=5) bcd_temp[3:0]=bcd_temp[3:0]+3;
    if(bcd_temp[7:4]>=5) bcd_temp[7:4]=bcd_temp[7:4]+3;
    if(bcd_temp[11:8]>=5) bcd_temp[11:8]=bcd_temp[11:8]+3;
    if(bcd_temp[15:12]>=5) bcd_temp[15:12]=bcd_temp[15:12]+3;
    bcd_temp={bcd_temp[14:0],bin[13-count]};
    count=count+1;
end
else
begin
    reset=1;
    bcd=bcd_temp;
end
endmodule
module DINO_DATA(clk_25M,dino_data,dino_adrs,title_adrs,obstacle_data,obstacle_adrs,title,score_adrs,score_t,go_adrs,game_over);
input clk_25M;
input [5:0] title_adrs,dino_adrs,go_adrs;
input [4:0] score_adrs;
input [6:0] obstacle_adrs;
reg count=0;
output reg [63:0] dino_data;
output reg [79:0] obstacle_data;
output reg [0:399] title;
output reg [0:99] score_t;
output reg [0:235] game_over;
always @(posedge clk_25M)
begin
    case(count)
    4'd0:
        begin
            case(dino_adrs)
                6'd00:dino_data<=64'b0000000000000000000000000000000000000000000000000000000000000000;
                6'd01:dino_data<=64'b0000001111111111111111111111100000000000000000000000000000000000;
                6'd02:dino_data<=64'b0000001111111111111111111111100000000000000000000000000000000000;
                6'd03:dino_data<=64'b0001111111111111111111111111111100000000000000000000000000000000;
                6'd04:dino_data<=64'b0001111111111111111111111111111100000000000000000000000000000000;
                6'd05:dino_data<=64'b0001111111111111111111100011111100000000000000000000000000000000;
                6'd06:dino_data<=64'b0001111111111111111111100011111100000000000000000000000000000000;
                6'd07:dino_data<=64'b0001111111111111111111100011111100000000000000000000000000000000;
                6'd08:dino_data<=64'b0001111111111111111111111111111100000000000000000000000000000000;
                6'd09:dino_data<=64'b0001111111111111111111111111111100000000000000000000000000000000;
                6'd10:dino_data<=64'b0001111111111111111111111111111100000000000000000000000000000000;
                6'd11:dino_data<=64'b0001111111111111111111111111111100000000000000000000000000000000;
                6'd12:dino_data<=64'b0001111111111111111111111111111100000000000000000000000000000000;
                6'd13:dino_data<=64'b0001111111111111111111111111111100000000000000000000000000000000;
                6'd14:dino_data<=64'b0001111111111111111111111111111100000000000000000000000000000000;
                6'd15:dino_data<=64'b0001111111111111111111111111111100000000000000000000000000000000;
                6'd16:dino_data<=64'b0000000000000000011111111111111100000000000000000000000000000000;
                6'd17:dino_data<=64'b0000000000000000001111111111111100000000000000000000000000000000;
                6'd18:dino_data<=64'b0000000000000000001111111111111100000000000000000000000000000000;
                6'd19:dino_data<=64'b0000000000000000011111111111111100000000000000000000000000000000;
                6'd20:dino_data<=64'b0000000001111111111111111111111100000000000000000000000000000000;
                6'd21:dino_data<=64'b0000000001111111111111111111111100000000000000000000000000000000;
                6'd22:dino_data<=64'b0000000000000000000011111111111110000000000000000000000000000000;
                6'd23:dino_data<=64'b0000000000000000000011111111111111100000000000000000000000011000;
                6'd24:dino_data<=64'b0000000000000000000011111111111111100000000000000000000000011000;
                6'd25:dino_data<=64'b0000000000000000000011111111111111110110000000000000000000011000;
                6'd26:dino_data<=64'b0000000000000000000011111111111111111110000000000000000000011000;
                6'd27:dino_data<=64'b0000000000000000000011111111111111111110000000000000000000011000;
                6'd28:dino_data<=64'b0000000000000001111111111111111111111111111100000000000011111000;
                6'd29:dino_data<=64'b0000000000000001111111111111111111111111111100000000000011111000;
                6'd30:dino_data<=64'b0000000000000001111111111111111111111111111100000000000011111000;
                6'd31:dino_data<=64'b0000000000000001100011111111111111111111111111100000011111111000;
                6'd32:dino_data<=64'b0000000000000001100011111111111111111111111111100000011111111000;
                6'd33:dino_data<=64'b0000000000000001100011111111111111111111111111100000011111111000;
                6'd34:dino_data<=64'b0000000000000000000011111111111111111111111111111111111111111000;
                6'd35:dino_data<=64'b0000000000000000000011111111111111111111111111111111111111111000;
                6'd36:dino_data<=64'b0000000000000000000011111111111111111111111111111111111111111000;
                6'd37:dino_data<=64'b0000000000000000000011111111111111111111111111111111111111111000;
                6'd38:dino_data<=64'b0000000000000000000011111111111111111111111111111111111111111000;
                6'd39:dino_data<=64'b0000000000000000000011111111111111111111111111111111111111100000;
                6'd40:dino_data<=64'b0000000000000000000011111111111111111111111111111111111111000000;
                6'd41:dino_data<=64'b0000000000000000000000011111111111111111111111111111111111000000;
                6'd42:dino_data<=64'b0000000000000000000000011111111111111111111111111111111100000000;
                6'd43:dino_data<=64'b0000000000000000000000011111111111111111111111111111111100000000;
                6'd44:dino_data<=64'b0000000000000000000000011111111111111111111111111111111000000000;
                6'd45:dino_data<=64'b0000000000000000000000011111111111111111111111111111111100000000;
                6'd46:dino_data<=64'b0000000000000000000000000011111111111111111111111111100000000000;
                6'd47:dino_data<=64'b0000000000000000000000000011111111111111111111111111100000000000;
                6'd48:dino_data<=64'b0000000000000000000000000011111111111111111111111111100000000000;
                6'd49:dino_data<=64'b0000000000000000000000000000011111111111111111111100000000000000;
                6'd50:dino_data<=64'b0000000000000000000000000000011111111111111111111100000000000000;
                6'd51:dino_data<=64'b0000000000000000000000000000011111111111111111111100000000000000;
                6'd52:dino_data<=64'b0000000000000000000000000000011111100001111111100000000000000000;
                6'd53:dino_data<=64'b0000000000000000000000000000011111100001111111100000000000000000;
                6'd54:dino_data<=64'b0000000000000000000000000000011111100001111111100000000000000000;
                6'd55:dino_data<=64'b0000000000000000000000000000011100000000001111100000000000000000;
                6'd56:dino_data<=64'b0000000000000000000000000000011100000000001111100000000000000000;
                6'd57:dino_data<=64'b0000000000000000000000000000011100000000001111100000000000000000;
                6'd58:dino_data<=64'b0000000000000000000000000000011100000000000011100000000000000000;
                6'd59:dino_data<=64'b0000000000000000000000000000011100000000000011100000000000000000;
                6'd60:dino_data<=64'b0000000000000000000000000000011100000000000011100000000000000000;
                6'd61:dino_data<=64'b0000000000000000000000000011111100000000001111100000000000000000;
                6'd62:dino_data<=64'b0000000000000000000000000011111100000000001111100000000000000000;
                6'd63:dino_data<=64'b0000000000000000000000000001011100000000001011100000000000000000;
            endcase
        end
    endcase
end
always @(posedge clk_25M)
begin
    case(obstacle_adrs)
        7'd00:obstacle_data<=60'b000000000000000000000000000000000000000000000000000000000000;
        7'd01:obstacle_data<=60'b000000000000000000000000000000000000000000000000000000000000;
        7'd02:obstacle_data<=60'b000000000000000000000000000000000000000000000000000000000000;
        7'd03:obstacle_data<=60'b000000000000000000000000000000000000000000000000000000000000;
        7'd04:obstacle_data<=60'b000000000000000000000000000000111111100000000000000000000000;
        7'd05:obstacle_data<=60'b000000000000000000000000000011111111110000000000000000000000;
        7'd06:obstacle_data<=60'b000000000000000000000000000111111111111000000000000000000000;
        7'd07:obstacle_data<=60'b000000000000000000000000000111111111111100000000000000000000;
        7'd08:obstacle_data<=60'b000000000000000000000000000111111111111100000000000000000000;
        7'd09:obstacle_data<=60'b000000000000000000000000001111111111111110000000000000000000;
        7'd10:obstacle_data<=60'b000000001110000000000000001111111111111110000000000000000000;
        7'd11:obstacle_data<=60'b000000011111000000000000001111111111111110000000000000000000;
        7'd12:obstacle_data<=60'b000000011111000000000000001111111111111110000000000000000000;
        7'd13:obstacle_data<=60'b000000111111100000000000011111111111111111000000000000000000;
        7'd14:obstacle_data<=60'b000000111111100000000000011111111111111111000000000000000000;
        7'd15:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd16:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd17:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd18:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd19:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd20:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd21:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd22:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd23:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd24:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd25:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd26:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd27:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd28:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd29:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd30:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd31:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd32:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd33:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd34:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd35:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd36:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd37:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd38:obstacle_data<=60'b000001111111110000000000011111111111111111000000000000000000;
        7'd39:obstacle_data<=60'b000001111111110000000000011111111111111111000000000001000000;
        7'd40:obstacle_data<=60'b000001111111110000000000011111111111111111000000001111110000;
        7'd41:obstacle_data<=60'b000001111111111000000000011111111111111111000000011111110000;
        7'd42:obstacle_data<=60'b000001111111111000000000011111111111111111000000011111111000;
        7'd43:obstacle_data<=60'b000001111111111000000000011111111111111111000000111111111000;
        7'd44:obstacle_data<=60'b000001111111111000000000011111111111111111000000111111111000;
        7'd45:obstacle_data<=60'b000001111111111100000000011111111111111111000001111111111000;
        7'd46:obstacle_data<=60'b000001111111111100000000011111111111111111000001111111111000;
        7'd47:obstacle_data<=60'b000001111111111100000000011111111111111111000011111111111000;
        7'd48:obstacle_data<=60'b000001111111111110000000011111111111111111000011111111111000;
        7'd49:obstacle_data<=60'b000001111111111111000000011111111111111111000011111111110000;
        7'd50:obstacle_data<=60'b000001111111111111000000011111111111111111000011111111110000;
        7'd51:obstacle_data<=60'b000000111111111111100000011111111111111111000111111111110000;
        7'd52:obstacle_data<=60'b000000011111111111111000011111111111111111000111111111100000;
        7'd53:obstacle_data<=60'b000000001111111111111100001111111111111111000111111111100000;
        7'd54:obstacle_data<=60'b000000000111111111111111001111111111111111001111111111000000;
        7'd55:obstacle_data<=60'b000000000011111111111111111111111111111111011111111111000000;
        7'd56:obstacle_data<=60'b000000000001111111111111111111111111111111111111111110000000;
        7'd57:obstacle_data<=60'b000000000000111111111111111111111111111111111111111100000000;
        7'd58:obstacle_data<=60'b000000000000001111111111111111111111111111111111111000000000;
        7'd59:obstacle_data<=60'b000000000000000011111111111111111111111111111111110000000000;
        7'd60:obstacle_data<=60'b000000000000000000001111111111111111111111111111000000000000;
        7'd61:obstacle_data<=60'b000000000000000000000000011111111111111111111100000000000000;
        7'd62:obstacle_data<=60'b000000000000000000000000001111111111111000000000000000000000;
        7'd63:obstacle_data<=60'b000000000000000000000000000111111111110000000000000000000000;
        7'd64:obstacle_data<=60'b000000000000000000000000000111111111110000000000000000000000;
        7'd65:obstacle_data<=60'b000000000000000000000000000111111111110000000000000000000000;
        7'd66:obstacle_data<=60'b000000000000000000000000000111111111110000000000000000000000;
        7'd67:obstacle_data<=60'b000000000000000000000000000111111111110000000000000000000000;
        7'd68:obstacle_data<=60'b000000000000000000000000000111111111110000000000000000000000;
        7'd69:obstacle_data<=60'b000000000000000000000000000111111111110000000000000000000000;
        7'd70:obstacle_data<=60'b000000000000000000000000000111111111110000000000000000000000;
        7'd71:obstacle_data<=60'b000000000000000000000000000011111111100000000000000000000000;
        7'd72:obstacle_data<=60'b000000000000000000000000000011111111100000000000000000000000;
        7'd73:obstacle_data<=60'b000000000000000000000000000011111111100000000000000000000000;
        7'd74:obstacle_data<=60'b000000000000000000000000000011111111100000000000000000000000;
        7'd75:obstacle_data<=60'b000000000000000000000000000011111111100000000000000000000000;
        7'd76:obstacle_data<=60'b000000000000000000000000001111111111111000000000000000000000;
        7'd77:obstacle_data<=60'b000000000000000000000000000000000000000000000000000000000000;
        7'd78:obstacle_data<=60'b000000000000000000000000000000000000000000000000000000000000;
        7'd79:obstacle_data<=60'b000000000000000000000000000000000000000000000000000000000000;
        default:
            obstacle_data<=obstacle_data;
    endcase
end
always @(posedge clk_25M)
begin
    case(title_adrs)
        6'd00:title<=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd01:title<=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd02:title<=400'b0001111111111111111111111111100000000000000000000011111111110000000001111111111000000000000000000011111111100000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000011111111111000000000000000000000001111111111111110000000000000000011111111111111000000000011111111111111111111111111111111111000;
        6'd03:title<=400'b0001111111111111111111111111111100000000000000000011111111110000000001111111111100000000000000000011111111100000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000011111111111000000000000000000000001111111111111110000000000000000111111111111111000000000011111111111111111111111111111111111000;
        6'd04:title<=400'b0001111111111111111111111111111110000000000000000011111111110000000001111111111100000000000000000011111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000111111111111100000000000000000000001111111111111111000000000000000111111111111111000000000011111111111111111111111111111111111000;
        6'd05:title<=400'b0001111111111111111111111111111111100000000000000011111111110000000001111111111110000000000000000011111111100000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000111111111111100000000000000000000001111111111111111000000000000000111111111111111000000000011111111111111111111111111111111111000;
        6'd06:title<=400'b0001111111111111111111111111111111110000000000000011111111110000000001111111111110000000000000000011111111100000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000001111111111111100000000000000000000001111111111111111000000000000000111111111111111000000000011111111111111111111111111111111111000;
        6'd07:title<=400'b0001111111111111111111111111111111111000000000000011111111110000000001111111111111000000000000000011111111100000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000000001111111111111110000000000000000000001111111111111111000000000000001111111111111111000000000011111111111111111111111111111111111000;
        6'd08:title<=400'b0001111111111111111111111111111111111100000000000011111111110000000001111111111111100000000000000011111111100000000000001111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000000001111111111111110000000000000000000001111111111111111100000000000001111111111111111000000000011111111111111111111111111111111111000;
        6'd09:title<=400'b0001111111111111111111111111111111111100000000000011111111110000000001111111111111100000000000000011111111100000000000001111111111111100000000111111111111111000000000000000000000000000000000000000000000000000001111111111111110000000111111111111111000000000000000000000011111111111111111000000000000000000001111111111111111100000000000001111111111111111000000000011111111111111111111111111111111111000;
        6'd10:title<=400'b0001111111110000000000000011111111111110000000000011111111110000000001111111111111110000000000000011111111100000000000011111111111110000000000001111111111111000000000000000000000000000000000000000000000000000011111111111110000000000000111111111111100000000000000000000011111111111111111000000000000000000001111111111111111100000000000001111111111111111000000000011111111100000000000000000000000000000;
        6'd11:title<=400'b0001111111110000000000000000111111111111000000000011111111110000000001111111111111111000000000000011111111100000000000111111111111000000000000000011111111111100000000000000000000000000000000000000000000000000011111111111100000000000000011111111111100000000000000000000111111111111111111000000000000000000001111111111111111100000000000011111111111111111000000000011111111100000000000000000000000000000;
        6'd12:title<=400'b0001111111110000000000000000011111111111000000000011111111110000000001111111111111111000000000000011111111100000000000111111111110000000000000000001111111111100000000000000000000000000000000000000000000000000111111111111000000000000000001111111111110000000000000000000111111111111111111100000000000000000001111111111111111110000000000011111111111111111000000000011111111100000000000000000000000000000;
        6'd13:title<=400'b0001111111110000000000000000001111111111000000000011111111110000000001111111111111111100000000000011111111100000000001111111111100000000000000000000111111111110000000000000000000000000000000000000000000000000111111111110000000000000000000111111111110000000000000000000111111111111111111100000000000000000001111111111111111110000000000011111111111111111000000000011111111100000000000000000000000000000;
        6'd14:title<=400'b0001111111110000000000000000001111111111100000000011111111110000000001111111111111111100000000000011111111100000000001111111111100000000000000000000011111111110000000000000000000000000000000000000000000000001111111111100000000000000000000011111111110000000000000000001111111111011111111110000000000000000001111111111111111110000000000011111111111111111000000000011111111100000000000000000000000000000;
        6'd15:title<=400'b0001111111110000000000000000000111111111100000000011111111110000000001111111111111111110000000000011111111100000000011111111111000000000000000000000011111111111000000000000000000000000000000000000000000000001111111111000000000000000000000011111110000000000000000000001111111110011111111110000000000000000001111111110111111111000000000111111111111111111000000000011111111100000000000000000000000000000;
        6'd16:title<=400'b0001111111110000000000000000000111111111100000000011111111110000000001111111111111111111000000000011111111100000000011111111110000000000000000000000001111111111000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110001111111110000000000000000001111111110111111111000000000111111110111111111000000000011111111100000000000000000000000000000;
        6'd17:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111111111111111000000000011111111100000000011111111110000000000000000000000001111111111000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000011111111110001111111111000000000000000001111111110011111111000000000111111110111111111000000000011111111100000000000000000000000000000;
        6'd18:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111111111111111100000000011111111100000000011111111110000000000000000000000001111111111000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000011111111100001111111111000000000000000001111111110011111111000000001111111110111111111000000000011111111100000000000000000000000000000;
        6'd19:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110111111111100000000011111111100000000011111111110000000000000000000000000111111111100000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000111111111100000111111111100000000000000001111111110011111111100000001111111110111111111000000000011111111110000000000000000000000000000;
        6'd20:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110111111111110000000011111111100000000111111111100000000000000000000000000111111111100000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000111111111000000111111111100000000000000001111111110011111111100000001111111100111111111000000000011111111111111111111111111111111100000;
        6'd21:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110011111111111000000011111111100000000111111111100000000000000000000000000111111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000111111111000000111111111100000000000000001111111110001111111100000001111111100111111111000000000011111111111111111111111111111111100000;
        6'd22:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110001111111111000000011111111100000000111111111100000000000000000000000000111111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000001111111111000000011111111110000000000000001111111110001111111100000011111111100111111111000000000011111111111111111111111111111111100000;
        6'd23:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110001111111111100000011111111100000000111111111100000000000000000000000000111111111100000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000001111111110000000011111111110000000000000001111111110001111111110000011111111000111111111000000000011111111111111111111111111111111100000;
        6'd24:title<=400'b0001111111110000000000000000000001111111110000000011111111110000000001111111110000011111111110000011111111100000000111111111100000000000000000000000000111111111100000000000000000000000000000000000000000000111111111100000000000000111111111111111111111000000000000011111111110000000001111111111000000000000001111111110000111111110000011111111000111111111000000000011111111111111111111111111111111100000;
        6'd25:title<=400'b0001111111110000000000000000000001111111110000000011111111110000000001111111110000011111111111000011111111100000000111111111100000000000000000000000000111111111100000000000000000000000000000000000000000000111111111100000000000000111111111111111111111000000000000011111111100000000001111111111000000000000001111111110000111111110000111111111000111111111000000000011111111111111111111111111111111100000;
        6'd26:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110000001111111111000011111111100000000111111111100000000000000000000000000111111111100000000000000000000000000000000000000000000111111111100000000000000111111111111111111111000000000000111111111100000000000111111111100000000000001111111110000111111111000111111110000111111111000000000011111111111111111111111111111111100000;
        6'd27:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110000001111111111100011111111100000000111111111100000000000000000000000000111111111100000000000000000000000000000000000000000000011111111100000000000000111111111111111111111000000000000111111111100000000000111111111100000000000001111111110000011111111000111111110000111111111000000000011111111110000000000000000000000000000;
        6'd28:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110000000111111111110011111111100000000111111111100000000000000000000000000111111111100000000000000000000000000000000000000000000011111111110000000000000111111111111111111111000000000001111111111000000000000111111111110000000000001111111110000011111111000111111110000111111111000000000011111111100000000000000000000000000000;
        6'd29:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110000000011111111110011111111100000000111111111100000000000000000000000000111111111100000000000000000000000000000000000000000000011111111110000000000000111111111111111111111000000000001111111111111111111111111111111110000000000001111111110000011111111101111111110000111111111000000000011111111100000000000000000000000000000;
        6'd30:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110000000011111111111011111111100000000011111111110000000000000000000000001111111111100000000000000000000000000000000000000000000011111111110000000000000111111111111111111111000000000001111111111111111111111111111111110000000000001111111110000011111111101111111100000111111111000000000011111111100000000000000000000000000000;
        6'd31:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110000000001111111111111111111100000000011111111110000000000000000000000001111111111000000000000000000000000000000000000000000000011111111110000000000000000000000001111111111000000000011111111111111111111111111111111111000000000001111111110000001111111101111111100000111111111000000000011111111100000000000000000000000000000;
        6'd32:title<=400'b0001111111110000000000000000000011111111110000000011111111110000000001111111110000000001111111111111111111100000000011111111110000000000000000000000001111111111000000000000000000000000000000000000000000000001111111111000000000000000000000001111111111000000000011111111111111111111111111111111111000000000001111111110000001111111111111111100000111111111000000000011111111100000000000000000000000000000;
        6'd33:title<=400'b0001111111110000000000000000000111111111100000000011111111110000000001111111110000000000111111111111111111100000000011111111111000000000000000000000011111111111000000000000000000000000000000000000000000000001111111111000000000000000000000001111111111000000000011111111111111111111111111111111111100000000001111111110000001111111111111111100000111111111000000000011111111100000000000000000000000000000;
        6'd34:title<=400'b0001111111110000000000000000000111111111100000000011111111110000000001111111110000000000011111111111111111100000000001111111111000000000000000000000011111111111000000000000000000000000000000000000000000000001111111111100000000000000000000001111111111000000000111111111111111111111111111111111111100000000001111111110000001111111111111111000000111111111000000000011111111100000000000000000000000000000;
        6'd35:title<=400'b0001111111110000000000000000000111111111100000000011111111110000000001111111110000000000011111111111111111100000000001111111111100000000000000000000111111111110000000000000000000000000000000000000000000000000111111111100000000000000000000001111111111000000000111111111111111111111111111111111111100000000001111111110000000111111111111111000000111111111000000000011111111100000000000000000000000000000;
        6'd36:title<=400'b0001111111110000000000000000001111111111000000000011111111110000000001111111110000000000001111111111111111100000000001111111111110000000000000000000111111111110000000000000000000000000000000000000000000000000111111111110000000000000000000001111111111000000001111111111111111111111111111111111111110000000001111111110000000111111111111111000000111111111000000000011111111100000000000000000000000000000;
        6'd37:title<=400'b0001111111110000000000000000011111111111000000000011111111110000000001111111110000000000000111111111111111100000000000111111111111000000000000000001111111111100000000000000000000000000000000000000000000000000011111111111000000000000000000011111111111000000001111111111000000000000000000011111111110000000001111111110000000111111111111111000000111111111000000000011111111100000000000000000000000000000;
        6'd38:title<=400'b0001111111110000000000000000111111111110000000000011111111110000000001111111110000000000000111111111111111100000000000111111111111100000000000000111111111111100000000000000000000000000000000000000000000000000011111111111100000000000000001111111111111000000001111111111000000000000000000011111111111000000001111111110000000111111111111110000000111111111000000000011111111100000000000000000000000000000;
        6'd39:title<=400'b0001111111110000000000000011111111111110000000000011111111110000000001111111110000000000000011111111111111100000000000011111111111111000000000001111111111111000000000000000000000000000000000000000000000000000001111111111111000000000000111111111111111000000011111111110000000000000000000001111111111000000001111111110000000011111111111110000000111111111000000000011111111110000000000000000000000000000;
        6'd40:title<=400'b0001111111111111111111111111111111111100000000000011111111110000000001111111110000000000000011111111111111100000000000001111111111111111000001111111111111110000000000000000000000000000000000000000000000000000001111111111111111000001111111111111111111000000011111111110000000000000000000001111111111000000001111111110000000011111111111110000000111111111000000000011111111111111111111111111111111111000;
        6'd41:title<=400'b0001111111111111111111111111111111111100000000000011111111110000000001111111110000000000000001111111111111100000000000001111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000111111111100000000000000000000001111111111100000001111111110000000011111111111110000000111111111000000000011111111111111111111111111111111111000;
        6'd42:title<=400'b0001111111111111111111111111111111111000000000000011111111110000000001111111110000000000000000111111111111100000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111110000000111111111100000000000000000000000111111111100000001111111110000000011111111111100000000111111111000000000011111111111111111111111111111111111000;
        6'd43:title<=400'b0001111111111111111111111111111111110000000000000011111111110000000001111111110000000000000000111111111111100000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111000000000111111111100000000000000000000000111111111110000001111111110000000001111111111100000000111111111000000000011111111111111111111111111111111111000;
        6'd44:title<=400'b0001111111111111111111111111111111000000000000000011111111110000000001111111110000000000000000011111111111100000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000001111111111000000000000000000000000011111111110000001111111110000000001111111111100000000111111111000000000011111111111111111111111111111111111000;
        6'd45:title<=400'b0001111111111111111111111111111110000000000000000011111111110000000001111111110000000000000000001111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111111000000000000000000000000011111111110000001111111110000000001111111111100000000111111111000000000011111111111111111111111111111111111000;
        6'd46:title<=400'b0001111111111111111111111111111000000000000000000011111111110000000001111111110000000000000000001111111111100000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000011111111111000000000000000000000000011111111111000001111111110000000001111111111000000000111111111000000000011111111111111111111111111111111111000;
        6'd47:title<=400'b0001111111111111111111111111000000000000000000000011111111110000000001111111110000000000000000000111111111100000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000011111111110000000000000000000000000001111111111000001111111110000000000111111111000000000111111111000000000011111111111111111111111111111111111000;
        6'd48:title<=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd49:title<=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
end
always @(posedge clk_25M)
begin
    case(score_adrs)
        5'd00:score_t<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd01:score_t<=100'b0000000110000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000;
        5'd02:score_t<=100'b0000111111110000000000011111110000000000011111111100000000001111111110000000001111111111110000000000;
        5'd03:score_t<=100'b0001111111111000000001111111111100000000111111111110000000001111111111100000001111111111110000000000;
        5'd04:score_t<=100'b0011111111111000000011111111111110000001111111111111000000001111111111110000001111111111110000000000;
        5'd05:score_t<=100'b0011100000011000000011110000011110000011110000001111100000001110000011110000001111000000000000000000;
        5'd06:score_t<=100'b0111100000000000000111100000000110000111100000000011100000001110000001111000001110000000000000000000;
        5'd07:score_t<=100'b0111000000000000000111000000000000000111000000000011110000001110000001111000001110000000000000000000;
        5'd08:score_t<=100'b0111000000000000001111000000000000000111000000000001110000001110000000111000001110000000000000000000;
        5'd09:score_t<=100'b0111000000000000001110000000000000001111000000000001110000001110000000111000001110000000000000000000;
        5'd10:score_t<=100'b0111100000000000001110000000000000001110000000000001111000001110000000111000001110000000000000001100;
        5'd11:score_t<=100'b0111100000000000011110000000000000001110000000000000111000001110000000111000001110000000000000001110;
        5'd12:score_t<=100'b0011110000000000011100000000000000001110000000000000111000001110000001111000001110000000000000001110;
        5'd13:score_t<=100'b0011111000000000011100000000000000001110000000000000111000001110000001110000001110000000000000001110;
        5'd14:score_t<=100'b0001111110000000011100000000000000001110000000000000111000001110000111100000001111111111100000001110;
        5'd15:score_t<=100'b0000111111000000011100000000000000001110000000000000111000001111111111100000001111111111100000000000;
        5'd16:score_t<=100'b0000011111110000011100000000000000011110000000000000111000001111111110000000001111111111100000000000;
        5'd17:score_t<=100'b0000000111111000011100000000000000001110000000000000111000001111111111000000001111000000000000000000;
        5'd18:score_t<=100'b0000000011111000011100000000000000001110000000000000111000001110000111000000001110000000000000000000;
        5'd19:score_t<=100'b0000000000111100011100000000000000001110000000000000111000001110000011100000001110000000000000000000;
        5'd20:score_t<=100'b0000000000111100011100000000000000001110000000000000111000001110000011100000001110000000000000000000;
        5'd21:score_t<=100'b0000000000011100011110000000000000001110000000000001111000001110000001110000001110000000000000000000;
        5'd22:score_t<=100'b0000000000011100001110000000000000001110000000000001110000001110000001110000001110000000000000000000;
        5'd23:score_t<=100'b0000000000011100001110000000000000001111000000000001110000001110000001110000001110000000000000000000;
        5'd24:score_t<=100'b0000000000011100001111000000000000000111000000000011110000001110000001111000001110000000000000000000;
        5'd25:score_t<=100'b0000000000011100000111000000000010000111100000000011100000001110000000111000001110000000000000000000;
        5'd26:score_t<=100'b0110000000111000000111100000001110000111100000000111100000001110000000111000001110000000000000001110;
        5'd27:score_t<=100'b0111100001111000000011111000111110000011111000011111000000001110000000111100001111000000000000001110;
        5'd28:score_t<=100'b0111111111110000000011111111111100000001111111111110000000001110000000011100001111111111111000001110;
        5'd29:score_t<=100'b0011111111100000000001111111111000000000111111111100000000001110000000011100001111111111111000001110;
        5'd30:score_t<=100'b0001111111000000000000011111100000000000001111111000000000001110000000011100000111111111111000001110;
        5'd31:score_t<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
end
always @(posedge clk_25M)
begin
    case(go_adrs)
        6'd00:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd01:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd02:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd03:game_over<=236'b00000000011111111111100000000000000000001111000000000000001111110000000000000000111110000001111111111111111111100000000000000000000000011111111110000000000111100000000000000000011110001111111111111111111100000011111111111111111100000000;
6'd04:game_over<=236'b00000001111111111111111000000000000000011111100000000000001111110000000000000001111110000001111111111111111111100000000000000000000001111111111111100000000011110000000000000000111100001111111111111111111100000011111111111111111111000000;
6'd05:game_over<=236'b00000011111111111111111100000000000000011111100000000000001111111000000000000001111110000001111111111111111111100000000000000000000111111111111111111000000011110000000000000000111100001111111111111111111100000011111111111111111111100000;
6'd06:game_over<=236'b00000111111000000001111110000000000000011111100000000000001111111000000000000001111110000001111000000000000000000000000000000000001111110000000011111100000001111000000000000000111000001111000000000000000000000011110000000000001111100000;
6'd07:game_over<=236'b00001111100000000000011110000000000000111111110000000000001111111000000000000011111110000001111000000000000000000000000000000000011111000000000000111100000001111000000000000001111000001111000000000000000000000011110000000000000111110000;
6'd08:game_over<=236'b00011111000000000000001111000000000000111001110000000000001111111100000000000011111110000001111000000000000000000000000000000000011110000000000000011110000001111000000000000001111000001111000000000000000000000011110000000000000011110000;
6'd09:game_over<=236'b00011110000000000000001111000000000000111001111000000000001111111100000000000011111110000001111000000000000000000000000000000000111100000000000000011111000000111100000000000001110000001111000000000000000000000011110000000000000001110000;
6'd10:game_over<=236'b00111100000000000000000111000000000001111001111000000000001111011100000000000111011110000001111000000000000000000000000000000000111100000000000000001111000000111100000000000011110000001111000000000000000000000011110000000000000001110000;
6'd11:game_over<=236'b00111100000000000000000100000000000001110000111100000000001111011110000000000111011110000001111000000000000000000000000000000001111000000000000000000111000000011100000000000011100000001111000000000000000000000011110000000000000001110000;
6'd12:game_over<=236'b00111100000000000000000000000000000011110000111100000000001111001110000000000111011110000001111000000000000000000000000000000001111000000000000000000111100000011110000000000111100000001111000000000000000000000011110000000000000011110000;
6'd13:game_over<=236'b01111000000000000000000000000000000011110000011100000000001111001110000000001110011110000001111000000000000000000000000000000001111000000000000000000111100000011110000000000111100000001111000000000000000000000011110000000000000011110000;
6'd14:game_over<=236'b01111000000000000000000000000000000011100000011110000000001111001111000000001110011110000001111000000000000000000000000000000001111000000000000000000111100000001110000000000111000000001111000000000000000000000011110000000000001111100000;
6'd15:game_over<=236'b01111000000000000000000000000000000111100000011110000000001111000111000000001110011110000001111111111111111111000000000000000001111000000000000000000111100000001111000000001111000000001111111111111111111000000011111111111111111111100000;
6'd16:game_over<=236'b01111000000000000000000000000000000111000000001111000000001111000111000000011100011110000001111111111111111111000000000000000001110000000000000000000111100000001111000000001111000000001111111111111111111000000011111111111111111110000000;
6'd17:game_over<=236'b01111000000000011111111111100000001111000000001111000000001111000111100000011100011110000001111111111111111111000000000000000001110000000000000000000111100000000111000000001110000000001111111111111111111000000011111111111111111000000000;
6'd18:game_over<=236'b01111000000000011111111111100000001111000000001111000000001111000011100000011100011110000001111000000000000000000000000000000001111000000000000000000111100000000111100000011110000000001111000000000000000000000011111111111111110000000000;
6'd19:game_over<=236'b01111000000000011111111111100000001111111111111111100000001111000011100000111000011110000001111000000000000000000000000000000001111000000000000000000111100000000011100000011100000000001111000000000000000000000011110000000011111000000000;
6'd20:game_over<=236'b01111000000000000000000111100000011111111111111111100000001111000011110000111000011110000001111000000000000000000000000000000001111000000000000000000111100000000011110000011100000000001111000000000000000000000011110000000001111100000000;
6'd21:game_over<=236'b00111100000000000000000111100000011111111111111111110000001111000001110000111000011110000001111000000000000000000000000000000001111000000000000000000111100000000011110000111100000000001111000000000000000000000011110000000000111110000000;
6'd22:game_over<=236'b00111100000000000000000111100000011110000000000011110000001111000001110001110000011110000001111000000000000000000000000000000000111000000000000000000111000000000001110000111000000000001111000000000000000000000011110000000000011110000000;
6'd23:game_over<=236'b00111100000000000000000111100000111100000000000011110000001111000001111001110000011110000001111000000000000000000000000000000000111100000000000000001111000000000001111001111000000000001111000000000000000000000011110000000000011111000000;
6'd24:game_over<=236'b00011110000000000000000111100000111100000000000001111000001111000000111001110000011110000001111000000000000000000000000000000000111110000000000000011111000000000000111001110000000000001111000000000000000000000011110000000000001111100000;
6'd25:game_over<=236'b00011111000000000000000111100001111000000000000001111000001111000000111011100000011110000001111000000000000000000000000000000000011110000000000000011110000000000000111001110000000000001111000000000000000000000011110000000000000111100000;
6'd26:game_over<=236'b00001111100000000000011111100001111000000000000000111100001111000000111111100000011110000001111000000000000000000000000000000000001111100000000001111100000000000000111111110000000000001111000000000000000000000011110000000000000111110000;
6'd27:game_over<=236'b00000111111100000001111111000001110000000000000000111100001111000000011111000000011110000001111000000000000000000000000000000000000111110000000011111100000000000000011111100000000000001111000000000000000000000011110000000000000011111000;
6'd28:game_over<=236'b00000011111111111111111110000011110000000000000000111110001111000000011111000000011110000001111111111111111111110000000000000000000011111111111111110000000000000000011111100000000000001111111111111111111110000011110000000000000001111000;
6'd29:game_over<=236'b00000000111111111111111000000011110000000000000000011110001111000000011111000000011110000001111111111111111111110000000000000000000001111111111111100000000000000000001111000000000000001111111111111111111110000011110000000000000001111100;
6'd30:game_over<=236'b00000000001111111111100000000011100000000000000000011110001111000000001110000000011110000001111111111111111111110000000000000000000000011111111110000000000000000000001111000000000000001111111111111111111110000011110000000000000000111100;
6'd31:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd32:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd33:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd34:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd35:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd36:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd37:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd38:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd39:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd40:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd41:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd42:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd43:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110111000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd44:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110111000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd45:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd46:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd47:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd48:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd49:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd50:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd51:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd52:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd53:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd54:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd55:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd56:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd57:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd58:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd59:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd60:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd61:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd62:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
6'd63:game_over<=236'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
end
endmodule

module SCORE_DATA(clk_25MHz,count,data,data_adrs);
input clk_25MHz;
input [4:0] data_adrs;
input [3:0] count;
output reg [0:19] data;
always @(posedge clk_25MHz)
begin
    case(count)
    4'd0:
        begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000011000000000;
        5'd03:data<=20'b00000011111111000000;
        5'd04:data<=20'b00000111111111100000;
        5'd05:data<=20'b00001111111111110000;
        5'd06:data<=20'b00001111111111110000;
        5'd07:data<=20'b00011111000011111000;
        5'd08:data<=20'b00011110000011111000;
        5'd09:data<=20'b00011110000001111000;
        5'd10:data<=20'b00111110000001111000;
        5'd11:data<=20'b00111110000001111000;
        5'd12:data<=20'b00111110000001111100;
        5'd13:data<=20'b00111100000001111100;
        5'd14:data<=20'b00111100000001111100;
        5'd15:data<=20'b00111100000001111100;
        5'd16:data<=20'b00111100000001111100;
        5'd17:data<=20'b00111100000001111100;
        5'd18:data<=20'b00111100000001111100;
        5'd19:data<=20'b00111110000001111100;
        5'd20:data<=20'b00111110000001111000;
        5'd21:data<=20'b00111110000001111000;
        5'd22:data<=20'b00111110000001111000;
        5'd23:data<=20'b00111110000011111000;
        5'd24:data<=20'b00011111000011111000;
        5'd25:data<=20'b00011111100111110000;
        5'd26:data<=20'b00011111111111110000;
        5'd27:data<=20'b00001111111111100000;
        5'd28:data<=20'b00000111111111000000;
        5'd29:data<=20'b00000011111110000000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;    
        endcase
        end
    4'd1:begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000000000000000;
        5'd04:data<=20'b00000001111000000000;
        5'd05:data<=20'b00000011111000000000;
        5'd06:data<=20'b00000111111000000000;
        5'd07:data<=20'b00011111111000000000;
        5'd08:data<=20'b00011111111000000000;
        5'd09:data<=20'b00011101111000000000;
        5'd10:data<=20'b00011001111000000000;
        5'd11:data<=20'b00000001111000000000;
        5'd12:data<=20'b00000001111000000000;
        5'd13:data<=20'b00000001111000000000;
        5'd14:data<=20'b00000001111000000000;
        5'd15:data<=20'b00000001111000000000;
        5'd16:data<=20'b00000001111000000000;
        5'd17:data<=20'b00000001111000000000;
        5'd18:data<=20'b00000001111000000000;
        5'd19:data<=20'b00000001111000000000;
        5'd20:data<=20'b00000001111000000000;
        5'd21:data<=20'b00000001111000000000;
        5'd22:data<=20'b00000001111000000000;
        5'd23:data<=20'b00000001111000000000;
        5'd24:data<=20'b00000001111000000000;
        5'd25:data<=20'b00000001111100000000;
        5'd26:data<=20'b00011111111111100000;
        5'd27:data<=20'b00011111111111100000;
        5'd28:data<=20'b00011111111111100000;
        5'd29:data<=20'b00011111111111100000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
        end
    4'd2:
        begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000001111100000000;
        5'd03:data<=20'b00000111111111000000;
        5'd04:data<=20'b00011111111111100000;
        5'd05:data<=20'b00011111111111100000;
        5'd06:data<=20'b00011111111111110000;
        5'd07:data<=20'b00011100011111110000;
        5'd08:data<=20'b00011000001111110000;
        5'd09:data<=20'b00000000000111110000;
        5'd10:data<=20'b00000000000111110000;
        5'd11:data<=20'b00000000000111110000;
        5'd12:data<=20'b00000000000111110000;
        5'd13:data<=20'b00000000001111110000;
        5'd14:data<=20'b00000000001111100000;
        5'd15:data<=20'b00000000001111100000;
        5'd16:data<=20'b00000000011111000000;
        5'd17:data<=20'b00000000111111000000;
        5'd18:data<=20'b00000000111110000000;
        5'd19:data<=20'b00000001111100000000;
        5'd20:data<=20'b00000011111000000000;
        5'd21:data<=20'b00000111111000000000;
        5'd22:data<=20'b00001111110000000000;
        5'd23:data<=20'b00001111100000000000;
        5'd24:data<=20'b00011111000000000000;
        5'd25:data<=20'b00011111111111111000;
        5'd26:data<=20'b00111111111111111000;
        5'd27:data<=20'b00111111111111111000;
        5'd28:data<=20'b00011111111111111000;
        5'd29:data<=20'b00011111111111110000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
        end
    4'd3:
        begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000011000000000;
            5'd03:data<=20'b00000111111111000000;
            5'd04:data<=20'b00001111111111100000;
            5'd05:data<=20'b00011111111111100000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011100001111110000;
            5'd08:data<=20'b00010000000111110000;
            5'd09:data<=20'b00000000000111110000;
            5'd10:data<=20'b00000000000111110000;
            5'd11:data<=20'b00000000000111110000;
            5'd12:data<=20'b00000000000111110000;
            5'd13:data<=20'b00000000001111100000;
            5'd14:data<=20'b00000111111111000000;
            5'd15:data<=20'b00001111111110000000;
            5'd16:data<=20'b00001111111111000000;
            5'd17:data<=20'b00000111111111110000;
            5'd18:data<=20'b00000000011111110000;
            5'd19:data<=20'b00000000000111111000;
            5'd20:data<=20'b00000000000011111000;
            5'd21:data<=20'b00000000000011111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011111000;
            5'd24:data<=20'b00010000000111111000;
            5'd25:data<=20'b00111100001111111000;
            5'd26:data<=20'b00111111111111110000;
            5'd27:data<=20'b00111111111111100000;
            5'd28:data<=20'b00011111111111000000;
            5'd29:data<=20'b00001111111110000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
            endcase
        end
    4'd4:
    begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000011111100000;
        5'd04:data<=20'b00000000011111100000;
        5'd05:data<=20'b00000000111111100000;
        5'd06:data<=20'b00000000111111100000;
        5'd07:data<=20'b00000001111111100000;
        5'd08:data<=20'b00000001111111100000;
        5'd09:data<=20'b00000011110111100000;
        5'd10:data<=20'b00000011110111100000;
        5'd11:data<=20'b00000111100111100000;
        5'd12:data<=20'b00000111100111100000;
        5'd13:data<=20'b00001111000111100000;
        5'd14:data<=20'b00001111000111100000;
        5'd15:data<=20'b00011110000111100000;
        5'd16:data<=20'b00011110000111100000;
        5'd17:data<=20'b00111100000111100000;
        5'd18:data<=20'b00111100000111100000;
        5'd19:data<=20'b00111000000111100000;
        5'd20:data<=20'b00111111111111111100;
        5'd21:data<=20'b00111111111111111100;
        5'd22:data<=20'b00111111111111111100;
        5'd23:data<=20'b00111111111111111100;
        5'd24:data<=20'b00000000000111110000;
        5'd25:data<=20'b00000000000111100000;
        5'd26:data<=20'b00000000000111100000;
        5'd27:data<=20'b00000000000111100000;
        5'd28:data<=20'b00000000000111100000;
        5'd29:data<=20'b00000000000111100000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd5:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00001111111111100000;
            5'd04:data<=20'b00011111111111110000;
            5'd05:data<=20'b00011111111111110000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011111111111100000;
            5'd08:data<=20'b00011110000000000000;
            5'd09:data<=20'b00011110000000000000;
            5'd10:data<=20'b00011110000000000000;
            5'd11:data<=20'b00011110000000000000;
            5'd12:data<=20'b00011110000000000000;
            5'd13:data<=20'b00011111111100000000;
            5'd14:data<=20'b00011111111111000000;
            5'd15:data<=20'b00011111111111100000;
            5'd16:data<=20'b00011111111111110000;
            5'd17:data<=20'b00001100011111111000;
            5'd18:data<=20'b00000000000111111000;
            5'd19:data<=20'b00000000000011111000;
            5'd20:data<=20'b00000000000011111000;
            5'd21:data<=20'b00000000000011111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011111000;
            5'd24:data<=20'b00000000000111111000;
            5'd25:data<=20'b00011000001111110000;
            5'd26:data<=20'b00011111111111110000;
            5'd27:data<=20'b00011111111111100000;
            5'd28:data<=20'b00011111111111000000;
            5'd29:data<=20'b00001111111100000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd6:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00000000111111110000;
            5'd04:data<=20'b00000011111111110000;
            5'd05:data<=20'b00000011111111110000;
            5'd06:data<=20'b00000111111111110000;
            5'd07:data<=20'b00001111100000000000;
            5'd08:data<=20'b00001111000000000000;
            5'd09:data<=20'b00011111000000000000;
            5'd10:data<=20'b00011110000000000000;
            5'd11:data<=20'b00011110000000000000;
            5'd12:data<=20'b00011110000000000000;
            5'd13:data<=20'b00011110011111000000;
            5'd14:data<=20'b00011111111111110000;
            5'd15:data<=20'b00011111111111111000;
            5'd16:data<=20'b00111111111111111000;
            5'd17:data<=20'b00111111000011111100;
            5'd18:data<=20'b00111110000001111100;
            5'd19:data<=20'b00011110000001111100;
            5'd20:data<=20'b00011110000001111100;
            5'd21:data<=20'b00011110000001111100;
            5'd22:data<=20'b00011110000001111100;
            5'd23:data<=20'b00011110000001111100;
            5'd24:data<=20'b00011111000001111000;
            5'd25:data<=20'b00011111100011111000;
            5'd26:data<=20'b00001111111111111000;
            5'd27:data<=20'b00001111111111110000;
            5'd28:data<=20'b00000111111111100000;
            5'd29:data<=20'b00000001111110000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd7:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00011111111111111000;
            5'd04:data<=20'b00111111111111111000;
            5'd05:data<=20'b00111111111111111000;
            5'd06:data<=20'b00111111111111111000;
            5'd07:data<=20'b00011111111111111000;
            5'd08:data<=20'b00000000000011111000;
            5'd09:data<=20'b00000000000011111000;
            5'd10:data<=20'b00000000000111110000;
            5'd11:data<=20'b00000000000111110000;
            5'd12:data<=20'b00000000000111110000;
            5'd13:data<=20'b00000000001111100000;
            5'd14:data<=20'b00000000001111100000;
            5'd15:data<=20'b00000000001111000000;
            5'd16:data<=20'b00000000011111000000;
            5'd17:data<=20'b00000000011111000000;
            5'd18:data<=20'b00000000111110000000;
            5'd19:data<=20'b00000000111110000000;
            5'd20:data<=20'b00000000111110000000;
            5'd21:data<=20'b00000001111100000000;
            5'd22:data<=20'b00000001111100000000;
            5'd23:data<=20'b00000011111100000000;
            5'd24:data<=20'b00000011111000000000;
            5'd25:data<=20'b00000011111000000000;
            5'd26:data<=20'b00000111110000000000;
            5'd27:data<=20'b00000111110000000000;
            5'd28:data<=20'b00000111110000000000;
            5'd29:data<=20'b00000111100000000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd8:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000001000000000;
            5'd03:data<=20'b00000011111111000000;
            5'd04:data<=20'b00000111111111100000;
            5'd05:data<=20'b00001111111111110000;
            5'd06:data<=20'b00011111101111111000;
            5'd07:data<=20'b00011111000011111000;
            5'd08:data<=20'b00011110000001111000;
            5'd09:data<=20'b00011110000001111000;
            5'd10:data<=20'b00011110000001111000;
            5'd11:data<=20'b00011111000011111000;
            5'd12:data<=20'b00011111000111110000;
            5'd13:data<=20'b00001111111111100000;
            5'd14:data<=20'b00001111111111100000;
            5'd15:data<=20'b00000111111111000000;
            5'd16:data<=20'b00000011111111000000;
            5'd17:data<=20'b00000111111111110000;
            5'd18:data<=20'b00001111101111110000;
            5'd19:data<=20'b00011111000111111000;
            5'd20:data<=20'b00011110000011111000;
            5'd21:data<=20'b00111110000001111100;
            5'd22:data<=20'b00111100000001111100;
            5'd23:data<=20'b00111100000001111100;
            5'd24:data<=20'b00111110000001111000;
            5'd25:data<=20'b00111111000011111000;
            5'd26:data<=20'b00011111111111111000;
            5'd27:data<=20'b00011111111111110000;
            5'd28:data<=20'b00001111111111100000;
            5'd29:data<=20'b00000011111111000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd9:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000011000000000;
            5'd03:data<=20'b00000011111111000000;
            5'd04:data<=20'b00000111111111100000;
            5'd05:data<=20'b00001111111111110000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011111000011111000;
            5'd08:data<=20'b00111110000011111000;
            5'd09:data<=20'b00111110000001111000;
            5'd10:data<=20'b00111100000001111000;
            5'd11:data<=20'b00111100000001111000;
            5'd12:data<=20'b00111110000001111000;
            5'd13:data<=20'b00111110000001111000;
            5'd14:data<=20'b00111110000001111000;
            5'd15:data<=20'b00011111000111111000;
            5'd16:data<=20'b00011111111111111000;
            5'd17:data<=20'b00011111111111111000;
            5'd18:data<=20'b00001111111111111000;
            5'd19:data<=20'b00000011111001111000;
            5'd20:data<=20'b00000000000001111000;
            5'd21:data<=20'b00000000000001111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011110000;
            5'd24:data<=20'b00000000000111110000;
            5'd25:data<=20'b00011000001111100000;
            5'd26:data<=20'b00011111111111100000;
            5'd27:data<=20'b00011111111111000000;
            5'd28:data<=20'b00011111111110000000;
            5'd29:data<=20'b00001111111000000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd10:
    begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000000000000000;
        5'd04:data<=20'b00000000000000000000;
        5'd05:data<=20'b00000000000000000000;
        5'd06:data<=20'b00000000000000000000;
        5'd07:data<=20'b00000000000000000000;
        5'd08:data<=20'b00000000000000000000;
        5'd09:data<=20'b00000000000000000000;
        5'd10:data<=20'b00000000011111000000;
        5'd11:data<=20'b00000000011111000000;
        5'd12:data<=20'b00000000011111000000;
        5'd13:data<=20'b00000000011111000000;
        5'd14:data<=20'b00000000000000000000;
        5'd15:data<=20'b00000000000000000000;
        5'd16:data<=20'b00000000000000000000;
        5'd17:data<=20'b00000000000000000000;
        5'd18:data<=20'b00000000000000000000;
        5'd19:data<=20'b00000000000000000000;
        5'd20:data<=20'b00000000000000000000;
        5'd21:data<=20'b00000000000000000000;
        5'd22:data<=20'b00000000000000000000;
        5'd23:data<=20'b00000000011111000000;
        5'd24:data<=20'b00000000011111000000;
        5'd25:data<=20'b00000000011111000000;
        5'd26:data<=20'b00000000011111000000;
        5'd27:data<=20'b00000000000000000000;
        5'd28:data<=20'b00000000000000000000;
        5'd29:data<=20'b00000000000000000000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
    end
    default:
        data<=0;    
    endcase
end
endmodule


